VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO Marmot
  CLASS BLOCK ;
  FOREIGN Marmot ;
  ORIGIN 0.000 0.000 ;
  SIZE 2880.000 BY 3480.000 ;
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 48.700 2884.800 49.900 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 2353.900 2884.800 2355.100 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 2584.420 2884.800 2585.620 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 2814.940 2884.800 2816.140 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 3045.460 2884.800 3046.660 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 3275.980 2884.800 3277.180 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2821.130 3479.000 2821.690 3484.800 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2502.350 3479.000 2502.910 3484.800 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2183.570 3479.000 2184.130 3484.800 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1864.790 3479.000 1865.350 3484.800 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1546.010 3479.000 1546.570 3484.800 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 279.220 2884.800 280.420 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1227.230 3479.000 1227.790 3484.800 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 908.450 3479.000 909.010 3484.800 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 589.670 3479.000 590.230 3484.800 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.890 3479.000 271.450 3484.800 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3426.260 1.000 3427.460 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3179.420 1.000 3180.620 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2932.580 1.000 2933.780 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2685.740 1.000 2686.940 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2438.900 1.000 2440.100 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2192.060 1.000 2193.260 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 509.740 2884.800 510.940 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1945.220 1.000 1946.420 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1698.380 1.000 1699.580 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1451.540 1.000 1452.740 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1204.700 1.000 1205.900 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 957.860 1.000 959.060 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 711.020 1.000 712.220 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 464.180 1.000 465.380 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 217.340 1.000 218.540 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 740.260 2884.800 741.460 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 970.780 2884.800 971.980 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 1201.300 2884.800 1202.500 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 1431.820 2884.800 1433.020 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 1662.340 2884.800 1663.540 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 1892.860 2884.800 1894.060 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 2123.380 2884.800 2124.580 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 202.380 2884.800 203.580 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 2507.580 2884.800 2508.780 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 2738.100 2884.800 2739.300 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 2968.620 2884.800 2969.820 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 3199.140 2884.800 3200.340 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 3429.660 2884.800 3430.860 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2608.610 3479.000 2609.170 3484.800 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2289.830 3479.000 2290.390 3484.800 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1971.050 3479.000 1971.610 3484.800 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1652.270 3479.000 1652.830 3484.800 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1333.490 3479.000 1334.050 3484.800 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 432.900 2884.800 434.100 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1014.710 3479.000 1015.270 3484.800 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 695.930 3479.000 696.490 3484.800 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 377.150 3479.000 377.710 3484.800 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.370 3479.000 58.930 3484.800 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3261.700 1.000 3262.900 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3014.860 1.000 3016.060 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2768.020 1.000 2769.220 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2521.180 1.000 2522.380 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2274.340 1.000 2275.540 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2027.500 1.000 2028.700 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 663.420 2884.800 664.620 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1780.660 1.000 1781.860 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1533.820 1.000 1535.020 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1286.980 1.000 1288.180 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1040.140 1.000 1041.340 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 793.300 1.000 794.500 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 546.460 1.000 547.660 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 299.620 1.000 300.820 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 52.780 1.000 53.980 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 893.940 2884.800 895.140 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 1124.460 2884.800 1125.660 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 1354.980 2884.800 1356.180 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 1585.500 2884.800 1586.700 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 1816.020 2884.800 1817.220 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 2046.540 2884.800 2047.740 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 2277.060 2884.800 2278.260 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 125.540 2884.800 126.740 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 2430.740 2884.800 2431.940 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 2661.260 2884.800 2662.460 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 2891.780 2884.800 2892.980 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 3122.300 2884.800 3123.500 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 3352.820 2884.800 3354.020 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2714.870 3479.000 2715.430 3484.800 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2396.090 3479.000 2396.650 3484.800 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2077.310 3479.000 2077.870 3484.800 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1758.530 3479.000 1759.090 3484.800 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1439.750 3479.000 1440.310 3484.800 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 356.060 2884.800 357.260 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1120.970 3479.000 1121.530 3484.800 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 802.190 3479.000 802.750 3484.800 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 483.410 3479.000 483.970 3484.800 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.630 3479.000 165.190 3484.800 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3343.980 1.000 3345.180 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3097.140 1.000 3098.340 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2850.300 1.000 2851.500 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2603.460 1.000 2604.660 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2356.620 1.000 2357.820 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2109.780 1.000 2110.980 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 586.580 2884.800 587.780 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1862.940 1.000 1864.140 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1616.100 1.000 1617.300 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1369.260 1.000 1370.460 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1122.420 1.000 1123.620 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 875.580 1.000 876.780 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 628.740 1.000 629.940 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 381.900 1.000 383.100 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 135.060 1.000 136.260 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 817.100 2884.800 818.300 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 1047.620 2884.800 1048.820 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 1278.140 2884.800 1279.340 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 1508.660 2884.800 1509.860 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 1739.180 2884.800 1740.380 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 1969.700 2884.800 1970.900 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 2200.220 2884.800 2201.420 ;
    END
  END io_out[9]
  PIN irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2786.630 -4.800 2787.190 1.000 ;
    END
  END irq[0]
  PIN irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2792.150 -4.800 2792.710 1.000 ;
    END
  END irq[1]
  PIN irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2797.670 -4.800 2798.230 1.000 ;
    END
  END irq[2]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 666.950 -4.800 667.510 1.000 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2322.950 -4.800 2323.510 1.000 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2339.510 -4.800 2340.070 1.000 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2356.070 -4.800 2356.630 1.000 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2372.630 -4.800 2373.190 1.000 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2389.190 -4.800 2389.750 1.000 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2405.750 -4.800 2406.310 1.000 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2422.310 -4.800 2422.870 1.000 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2438.870 -4.800 2439.430 1.000 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2455.430 -4.800 2455.990 1.000 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2471.990 -4.800 2472.550 1.000 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 832.550 -4.800 833.110 1.000 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2488.550 -4.800 2489.110 1.000 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2505.110 -4.800 2505.670 1.000 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2521.670 -4.800 2522.230 1.000 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2538.230 -4.800 2538.790 1.000 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2554.790 -4.800 2555.350 1.000 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2571.350 -4.800 2571.910 1.000 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2587.910 -4.800 2588.470 1.000 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2604.470 -4.800 2605.030 1.000 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2621.030 -4.800 2621.590 1.000 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2637.590 -4.800 2638.150 1.000 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 849.110 -4.800 849.670 1.000 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2654.150 -4.800 2654.710 1.000 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2670.710 -4.800 2671.270 1.000 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2687.270 -4.800 2687.830 1.000 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2703.830 -4.800 2704.390 1.000 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2720.390 -4.800 2720.950 1.000 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2736.950 -4.800 2737.510 1.000 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2753.510 -4.800 2754.070 1.000 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2770.070 -4.800 2770.630 1.000 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 865.670 -4.800 866.230 1.000 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 882.230 -4.800 882.790 1.000 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 898.790 -4.800 899.350 1.000 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 915.350 -4.800 915.910 1.000 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 931.910 -4.800 932.470 1.000 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 948.470 -4.800 949.030 1.000 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 965.030 -4.800 965.590 1.000 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 981.590 -4.800 982.150 1.000 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 683.510 -4.800 684.070 1.000 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 998.150 -4.800 998.710 1.000 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1014.710 -4.800 1015.270 1.000 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1031.270 -4.800 1031.830 1.000 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1047.830 -4.800 1048.390 1.000 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1064.390 -4.800 1064.950 1.000 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1080.950 -4.800 1081.510 1.000 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1097.510 -4.800 1098.070 1.000 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1114.070 -4.800 1114.630 1.000 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1130.630 -4.800 1131.190 1.000 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1147.190 -4.800 1147.750 1.000 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 700.070 -4.800 700.630 1.000 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1163.750 -4.800 1164.310 1.000 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1180.310 -4.800 1180.870 1.000 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1196.870 -4.800 1197.430 1.000 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1213.430 -4.800 1213.990 1.000 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1229.990 -4.800 1230.550 1.000 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1246.550 -4.800 1247.110 1.000 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1263.110 -4.800 1263.670 1.000 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1279.670 -4.800 1280.230 1.000 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1296.230 -4.800 1296.790 1.000 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1312.790 -4.800 1313.350 1.000 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 716.630 -4.800 717.190 1.000 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1329.350 -4.800 1329.910 1.000 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1345.910 -4.800 1346.470 1.000 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1362.470 -4.800 1363.030 1.000 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1379.030 -4.800 1379.590 1.000 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1395.590 -4.800 1396.150 1.000 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1412.150 -4.800 1412.710 1.000 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1428.710 -4.800 1429.270 1.000 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1445.270 -4.800 1445.830 1.000 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1461.830 -4.800 1462.390 1.000 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1478.390 -4.800 1478.950 1.000 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 733.190 -4.800 733.750 1.000 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1494.950 -4.800 1495.510 1.000 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1511.510 -4.800 1512.070 1.000 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1528.070 -4.800 1528.630 1.000 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1544.630 -4.800 1545.190 1.000 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1561.190 -4.800 1561.750 1.000 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1577.750 -4.800 1578.310 1.000 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1594.310 -4.800 1594.870 1.000 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1610.870 -4.800 1611.430 1.000 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1627.430 -4.800 1627.990 1.000 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1643.990 -4.800 1644.550 1.000 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 749.750 -4.800 750.310 1.000 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1660.550 -4.800 1661.110 1.000 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1677.110 -4.800 1677.670 1.000 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1693.670 -4.800 1694.230 1.000 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1710.230 -4.800 1710.790 1.000 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1726.790 -4.800 1727.350 1.000 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1743.350 -4.800 1743.910 1.000 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1759.910 -4.800 1760.470 1.000 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1776.470 -4.800 1777.030 1.000 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1793.030 -4.800 1793.590 1.000 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1809.590 -4.800 1810.150 1.000 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 766.310 -4.800 766.870 1.000 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1826.150 -4.800 1826.710 1.000 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1842.710 -4.800 1843.270 1.000 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1859.270 -4.800 1859.830 1.000 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1875.830 -4.800 1876.390 1.000 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1892.390 -4.800 1892.950 1.000 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1908.950 -4.800 1909.510 1.000 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1925.510 -4.800 1926.070 1.000 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1942.070 -4.800 1942.630 1.000 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1958.630 -4.800 1959.190 1.000 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1975.190 -4.800 1975.750 1.000 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 782.870 -4.800 783.430 1.000 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1991.750 -4.800 1992.310 1.000 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2008.310 -4.800 2008.870 1.000 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2024.870 -4.800 2025.430 1.000 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2041.430 -4.800 2041.990 1.000 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2057.990 -4.800 2058.550 1.000 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2074.550 -4.800 2075.110 1.000 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2091.110 -4.800 2091.670 1.000 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2107.670 -4.800 2108.230 1.000 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2124.230 -4.800 2124.790 1.000 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2140.790 -4.800 2141.350 1.000 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 799.430 -4.800 799.990 1.000 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2157.350 -4.800 2157.910 1.000 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2173.910 -4.800 2174.470 1.000 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2190.470 -4.800 2191.030 1.000 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2207.030 -4.800 2207.590 1.000 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2223.590 -4.800 2224.150 1.000 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2240.150 -4.800 2240.710 1.000 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2256.710 -4.800 2257.270 1.000 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2273.270 -4.800 2273.830 1.000 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2289.830 -4.800 2290.390 1.000 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2306.390 -4.800 2306.950 1.000 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 815.990 -4.800 816.550 1.000 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 672.470 -4.800 673.030 1.000 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2328.470 -4.800 2329.030 1.000 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2345.030 -4.800 2345.590 1.000 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2361.590 -4.800 2362.150 1.000 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2378.150 -4.800 2378.710 1.000 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2394.710 -4.800 2395.270 1.000 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2411.270 -4.800 2411.830 1.000 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2427.830 -4.800 2428.390 1.000 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2444.390 -4.800 2444.950 1.000 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2460.950 -4.800 2461.510 1.000 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2477.510 -4.800 2478.070 1.000 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 838.070 -4.800 838.630 1.000 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2494.070 -4.800 2494.630 1.000 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2510.630 -4.800 2511.190 1.000 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2527.190 -4.800 2527.750 1.000 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2543.750 -4.800 2544.310 1.000 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2560.310 -4.800 2560.870 1.000 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2576.870 -4.800 2577.430 1.000 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2593.430 -4.800 2593.990 1.000 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2609.990 -4.800 2610.550 1.000 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2626.550 -4.800 2627.110 1.000 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2643.110 -4.800 2643.670 1.000 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 854.630 -4.800 855.190 1.000 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2659.670 -4.800 2660.230 1.000 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2676.230 -4.800 2676.790 1.000 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2692.790 -4.800 2693.350 1.000 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2709.350 -4.800 2709.910 1.000 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2725.910 -4.800 2726.470 1.000 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2742.470 -4.800 2743.030 1.000 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2759.030 -4.800 2759.590 1.000 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2775.590 -4.800 2776.150 1.000 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 871.190 -4.800 871.750 1.000 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 887.750 -4.800 888.310 1.000 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 904.310 -4.800 904.870 1.000 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 920.870 -4.800 921.430 1.000 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 937.430 -4.800 937.990 1.000 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 953.990 -4.800 954.550 1.000 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 970.550 -4.800 971.110 1.000 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 987.110 -4.800 987.670 1.000 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 689.030 -4.800 689.590 1.000 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1003.670 -4.800 1004.230 1.000 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1020.230 -4.800 1020.790 1.000 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1036.790 -4.800 1037.350 1.000 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1053.350 -4.800 1053.910 1.000 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1069.910 -4.800 1070.470 1.000 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1086.470 -4.800 1087.030 1.000 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1103.030 -4.800 1103.590 1.000 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1119.590 -4.800 1120.150 1.000 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1136.150 -4.800 1136.710 1.000 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1152.710 -4.800 1153.270 1.000 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 705.590 -4.800 706.150 1.000 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1169.270 -4.800 1169.830 1.000 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1185.830 -4.800 1186.390 1.000 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1202.390 -4.800 1202.950 1.000 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1218.950 -4.800 1219.510 1.000 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1235.510 -4.800 1236.070 1.000 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1252.070 -4.800 1252.630 1.000 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1268.630 -4.800 1269.190 1.000 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1285.190 -4.800 1285.750 1.000 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1301.750 -4.800 1302.310 1.000 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1318.310 -4.800 1318.870 1.000 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 722.150 -4.800 722.710 1.000 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1334.870 -4.800 1335.430 1.000 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1351.430 -4.800 1351.990 1.000 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1367.990 -4.800 1368.550 1.000 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1384.550 -4.800 1385.110 1.000 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1401.110 -4.800 1401.670 1.000 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1417.670 -4.800 1418.230 1.000 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1434.230 -4.800 1434.790 1.000 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1450.790 -4.800 1451.350 1.000 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1467.350 -4.800 1467.910 1.000 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1483.910 -4.800 1484.470 1.000 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 738.710 -4.800 739.270 1.000 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1500.470 -4.800 1501.030 1.000 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1517.030 -4.800 1517.590 1.000 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1533.590 -4.800 1534.150 1.000 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1550.150 -4.800 1550.710 1.000 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1566.710 -4.800 1567.270 1.000 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1583.270 -4.800 1583.830 1.000 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1599.830 -4.800 1600.390 1.000 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1616.390 -4.800 1616.950 1.000 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1632.950 -4.800 1633.510 1.000 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1649.510 -4.800 1650.070 1.000 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 755.270 -4.800 755.830 1.000 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1666.070 -4.800 1666.630 1.000 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1682.630 -4.800 1683.190 1.000 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1699.190 -4.800 1699.750 1.000 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1715.750 -4.800 1716.310 1.000 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1732.310 -4.800 1732.870 1.000 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1748.870 -4.800 1749.430 1.000 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1765.430 -4.800 1765.990 1.000 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1781.990 -4.800 1782.550 1.000 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1798.550 -4.800 1799.110 1.000 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1815.110 -4.800 1815.670 1.000 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 771.830 -4.800 772.390 1.000 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1831.670 -4.800 1832.230 1.000 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1848.230 -4.800 1848.790 1.000 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1864.790 -4.800 1865.350 1.000 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1881.350 -4.800 1881.910 1.000 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1897.910 -4.800 1898.470 1.000 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1914.470 -4.800 1915.030 1.000 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1931.030 -4.800 1931.590 1.000 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1947.590 -4.800 1948.150 1.000 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1964.150 -4.800 1964.710 1.000 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1980.710 -4.800 1981.270 1.000 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 788.390 -4.800 788.950 1.000 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1997.270 -4.800 1997.830 1.000 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2013.830 -4.800 2014.390 1.000 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2030.390 -4.800 2030.950 1.000 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2046.950 -4.800 2047.510 1.000 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2063.510 -4.800 2064.070 1.000 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2080.070 -4.800 2080.630 1.000 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2096.630 -4.800 2097.190 1.000 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2113.190 -4.800 2113.750 1.000 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2129.750 -4.800 2130.310 1.000 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2146.310 -4.800 2146.870 1.000 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 804.950 -4.800 805.510 1.000 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2162.870 -4.800 2163.430 1.000 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2179.430 -4.800 2179.990 1.000 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2195.990 -4.800 2196.550 1.000 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2212.550 -4.800 2213.110 1.000 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2229.110 -4.800 2229.670 1.000 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2245.670 -4.800 2246.230 1.000 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2262.230 -4.800 2262.790 1.000 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2278.790 -4.800 2279.350 1.000 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2295.350 -4.800 2295.910 1.000 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2311.910 -4.800 2312.470 1.000 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 821.510 -4.800 822.070 1.000 ;
    END
  END la_data_out[9]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 677.990 -4.800 678.550 1.000 ;
    END
  END la_oenb[0]
  PIN la_oenb[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2333.990 -4.800 2334.550 1.000 ;
    END
  END la_oenb[100]
  PIN la_oenb[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2350.550 -4.800 2351.110 1.000 ;
    END
  END la_oenb[101]
  PIN la_oenb[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2367.110 -4.800 2367.670 1.000 ;
    END
  END la_oenb[102]
  PIN la_oenb[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2383.670 -4.800 2384.230 1.000 ;
    END
  END la_oenb[103]
  PIN la_oenb[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2400.230 -4.800 2400.790 1.000 ;
    END
  END la_oenb[104]
  PIN la_oenb[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2416.790 -4.800 2417.350 1.000 ;
    END
  END la_oenb[105]
  PIN la_oenb[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2433.350 -4.800 2433.910 1.000 ;
    END
  END la_oenb[106]
  PIN la_oenb[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2449.910 -4.800 2450.470 1.000 ;
    END
  END la_oenb[107]
  PIN la_oenb[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2466.470 -4.800 2467.030 1.000 ;
    END
  END la_oenb[108]
  PIN la_oenb[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2483.030 -4.800 2483.590 1.000 ;
    END
  END la_oenb[109]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 843.590 -4.800 844.150 1.000 ;
    END
  END la_oenb[10]
  PIN la_oenb[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2499.590 -4.800 2500.150 1.000 ;
    END
  END la_oenb[110]
  PIN la_oenb[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2516.150 -4.800 2516.710 1.000 ;
    END
  END la_oenb[111]
  PIN la_oenb[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2532.710 -4.800 2533.270 1.000 ;
    END
  END la_oenb[112]
  PIN la_oenb[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2549.270 -4.800 2549.830 1.000 ;
    END
  END la_oenb[113]
  PIN la_oenb[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2565.830 -4.800 2566.390 1.000 ;
    END
  END la_oenb[114]
  PIN la_oenb[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2582.390 -4.800 2582.950 1.000 ;
    END
  END la_oenb[115]
  PIN la_oenb[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2598.950 -4.800 2599.510 1.000 ;
    END
  END la_oenb[116]
  PIN la_oenb[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2615.510 -4.800 2616.070 1.000 ;
    END
  END la_oenb[117]
  PIN la_oenb[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2632.070 -4.800 2632.630 1.000 ;
    END
  END la_oenb[118]
  PIN la_oenb[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2648.630 -4.800 2649.190 1.000 ;
    END
  END la_oenb[119]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 860.150 -4.800 860.710 1.000 ;
    END
  END la_oenb[11]
  PIN la_oenb[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2665.190 -4.800 2665.750 1.000 ;
    END
  END la_oenb[120]
  PIN la_oenb[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2681.750 -4.800 2682.310 1.000 ;
    END
  END la_oenb[121]
  PIN la_oenb[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2698.310 -4.800 2698.870 1.000 ;
    END
  END la_oenb[122]
  PIN la_oenb[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2714.870 -4.800 2715.430 1.000 ;
    END
  END la_oenb[123]
  PIN la_oenb[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2731.430 -4.800 2731.990 1.000 ;
    END
  END la_oenb[124]
  PIN la_oenb[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2747.990 -4.800 2748.550 1.000 ;
    END
  END la_oenb[125]
  PIN la_oenb[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2764.550 -4.800 2765.110 1.000 ;
    END
  END la_oenb[126]
  PIN la_oenb[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2781.110 -4.800 2781.670 1.000 ;
    END
  END la_oenb[127]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 876.710 -4.800 877.270 1.000 ;
    END
  END la_oenb[12]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 893.270 -4.800 893.830 1.000 ;
    END
  END la_oenb[13]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 909.830 -4.800 910.390 1.000 ;
    END
  END la_oenb[14]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 926.390 -4.800 926.950 1.000 ;
    END
  END la_oenb[15]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 942.950 -4.800 943.510 1.000 ;
    END
  END la_oenb[16]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 959.510 -4.800 960.070 1.000 ;
    END
  END la_oenb[17]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 976.070 -4.800 976.630 1.000 ;
    END
  END la_oenb[18]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 992.630 -4.800 993.190 1.000 ;
    END
  END la_oenb[19]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 694.550 -4.800 695.110 1.000 ;
    END
  END la_oenb[1]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1009.190 -4.800 1009.750 1.000 ;
    END
  END la_oenb[20]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1025.750 -4.800 1026.310 1.000 ;
    END
  END la_oenb[21]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1042.310 -4.800 1042.870 1.000 ;
    END
  END la_oenb[22]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1058.870 -4.800 1059.430 1.000 ;
    END
  END la_oenb[23]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1075.430 -4.800 1075.990 1.000 ;
    END
  END la_oenb[24]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1091.990 -4.800 1092.550 1.000 ;
    END
  END la_oenb[25]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1108.550 -4.800 1109.110 1.000 ;
    END
  END la_oenb[26]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1125.110 -4.800 1125.670 1.000 ;
    END
  END la_oenb[27]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1141.670 -4.800 1142.230 1.000 ;
    END
  END la_oenb[28]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1158.230 -4.800 1158.790 1.000 ;
    END
  END la_oenb[29]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 711.110 -4.800 711.670 1.000 ;
    END
  END la_oenb[2]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1174.790 -4.800 1175.350 1.000 ;
    END
  END la_oenb[30]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1191.350 -4.800 1191.910 1.000 ;
    END
  END la_oenb[31]
  PIN la_oenb[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1207.910 -4.800 1208.470 1.000 ;
    END
  END la_oenb[32]
  PIN la_oenb[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1224.470 -4.800 1225.030 1.000 ;
    END
  END la_oenb[33]
  PIN la_oenb[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1241.030 -4.800 1241.590 1.000 ;
    END
  END la_oenb[34]
  PIN la_oenb[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1257.590 -4.800 1258.150 1.000 ;
    END
  END la_oenb[35]
  PIN la_oenb[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1274.150 -4.800 1274.710 1.000 ;
    END
  END la_oenb[36]
  PIN la_oenb[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1290.710 -4.800 1291.270 1.000 ;
    END
  END la_oenb[37]
  PIN la_oenb[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1307.270 -4.800 1307.830 1.000 ;
    END
  END la_oenb[38]
  PIN la_oenb[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1323.830 -4.800 1324.390 1.000 ;
    END
  END la_oenb[39]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 727.670 -4.800 728.230 1.000 ;
    END
  END la_oenb[3]
  PIN la_oenb[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1340.390 -4.800 1340.950 1.000 ;
    END
  END la_oenb[40]
  PIN la_oenb[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1356.950 -4.800 1357.510 1.000 ;
    END
  END la_oenb[41]
  PIN la_oenb[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1373.510 -4.800 1374.070 1.000 ;
    END
  END la_oenb[42]
  PIN la_oenb[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1390.070 -4.800 1390.630 1.000 ;
    END
  END la_oenb[43]
  PIN la_oenb[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1406.630 -4.800 1407.190 1.000 ;
    END
  END la_oenb[44]
  PIN la_oenb[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1423.190 -4.800 1423.750 1.000 ;
    END
  END la_oenb[45]
  PIN la_oenb[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1439.750 -4.800 1440.310 1.000 ;
    END
  END la_oenb[46]
  PIN la_oenb[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1456.310 -4.800 1456.870 1.000 ;
    END
  END la_oenb[47]
  PIN la_oenb[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1472.870 -4.800 1473.430 1.000 ;
    END
  END la_oenb[48]
  PIN la_oenb[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1489.430 -4.800 1489.990 1.000 ;
    END
  END la_oenb[49]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 744.230 -4.800 744.790 1.000 ;
    END
  END la_oenb[4]
  PIN la_oenb[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1505.990 -4.800 1506.550 1.000 ;
    END
  END la_oenb[50]
  PIN la_oenb[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1522.550 -4.800 1523.110 1.000 ;
    END
  END la_oenb[51]
  PIN la_oenb[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1539.110 -4.800 1539.670 1.000 ;
    END
  END la_oenb[52]
  PIN la_oenb[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1555.670 -4.800 1556.230 1.000 ;
    END
  END la_oenb[53]
  PIN la_oenb[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1572.230 -4.800 1572.790 1.000 ;
    END
  END la_oenb[54]
  PIN la_oenb[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1588.790 -4.800 1589.350 1.000 ;
    END
  END la_oenb[55]
  PIN la_oenb[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1605.350 -4.800 1605.910 1.000 ;
    END
  END la_oenb[56]
  PIN la_oenb[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1621.910 -4.800 1622.470 1.000 ;
    END
  END la_oenb[57]
  PIN la_oenb[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1638.470 -4.800 1639.030 1.000 ;
    END
  END la_oenb[58]
  PIN la_oenb[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1655.030 -4.800 1655.590 1.000 ;
    END
  END la_oenb[59]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 760.790 -4.800 761.350 1.000 ;
    END
  END la_oenb[5]
  PIN la_oenb[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1671.590 -4.800 1672.150 1.000 ;
    END
  END la_oenb[60]
  PIN la_oenb[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1688.150 -4.800 1688.710 1.000 ;
    END
  END la_oenb[61]
  PIN la_oenb[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1704.710 -4.800 1705.270 1.000 ;
    END
  END la_oenb[62]
  PIN la_oenb[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1721.270 -4.800 1721.830 1.000 ;
    END
  END la_oenb[63]
  PIN la_oenb[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1737.830 -4.800 1738.390 1.000 ;
    END
  END la_oenb[64]
  PIN la_oenb[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1754.390 -4.800 1754.950 1.000 ;
    END
  END la_oenb[65]
  PIN la_oenb[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1770.950 -4.800 1771.510 1.000 ;
    END
  END la_oenb[66]
  PIN la_oenb[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1787.510 -4.800 1788.070 1.000 ;
    END
  END la_oenb[67]
  PIN la_oenb[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1804.070 -4.800 1804.630 1.000 ;
    END
  END la_oenb[68]
  PIN la_oenb[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1820.630 -4.800 1821.190 1.000 ;
    END
  END la_oenb[69]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 777.350 -4.800 777.910 1.000 ;
    END
  END la_oenb[6]
  PIN la_oenb[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1837.190 -4.800 1837.750 1.000 ;
    END
  END la_oenb[70]
  PIN la_oenb[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1853.750 -4.800 1854.310 1.000 ;
    END
  END la_oenb[71]
  PIN la_oenb[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1870.310 -4.800 1870.870 1.000 ;
    END
  END la_oenb[72]
  PIN la_oenb[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1886.870 -4.800 1887.430 1.000 ;
    END
  END la_oenb[73]
  PIN la_oenb[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1903.430 -4.800 1903.990 1.000 ;
    END
  END la_oenb[74]
  PIN la_oenb[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1919.990 -4.800 1920.550 1.000 ;
    END
  END la_oenb[75]
  PIN la_oenb[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1936.550 -4.800 1937.110 1.000 ;
    END
  END la_oenb[76]
  PIN la_oenb[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1953.110 -4.800 1953.670 1.000 ;
    END
  END la_oenb[77]
  PIN la_oenb[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1969.670 -4.800 1970.230 1.000 ;
    END
  END la_oenb[78]
  PIN la_oenb[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1986.230 -4.800 1986.790 1.000 ;
    END
  END la_oenb[79]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 793.910 -4.800 794.470 1.000 ;
    END
  END la_oenb[7]
  PIN la_oenb[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2002.790 -4.800 2003.350 1.000 ;
    END
  END la_oenb[80]
  PIN la_oenb[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2019.350 -4.800 2019.910 1.000 ;
    END
  END la_oenb[81]
  PIN la_oenb[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2035.910 -4.800 2036.470 1.000 ;
    END
  END la_oenb[82]
  PIN la_oenb[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2052.470 -4.800 2053.030 1.000 ;
    END
  END la_oenb[83]
  PIN la_oenb[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2069.030 -4.800 2069.590 1.000 ;
    END
  END la_oenb[84]
  PIN la_oenb[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2085.590 -4.800 2086.150 1.000 ;
    END
  END la_oenb[85]
  PIN la_oenb[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2102.150 -4.800 2102.710 1.000 ;
    END
  END la_oenb[86]
  PIN la_oenb[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2118.710 -4.800 2119.270 1.000 ;
    END
  END la_oenb[87]
  PIN la_oenb[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2135.270 -4.800 2135.830 1.000 ;
    END
  END la_oenb[88]
  PIN la_oenb[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2151.830 -4.800 2152.390 1.000 ;
    END
  END la_oenb[89]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 810.470 -4.800 811.030 1.000 ;
    END
  END la_oenb[8]
  PIN la_oenb[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2168.390 -4.800 2168.950 1.000 ;
    END
  END la_oenb[90]
  PIN la_oenb[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2184.950 -4.800 2185.510 1.000 ;
    END
  END la_oenb[91]
  PIN la_oenb[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2201.510 -4.800 2202.070 1.000 ;
    END
  END la_oenb[92]
  PIN la_oenb[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2218.070 -4.800 2218.630 1.000 ;
    END
  END la_oenb[93]
  PIN la_oenb[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2234.630 -4.800 2235.190 1.000 ;
    END
  END la_oenb[94]
  PIN la_oenb[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2251.190 -4.800 2251.750 1.000 ;
    END
  END la_oenb[95]
  PIN la_oenb[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2267.750 -4.800 2268.310 1.000 ;
    END
  END la_oenb[96]
  PIN la_oenb[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2284.310 -4.800 2284.870 1.000 ;
    END
  END la_oenb[97]
  PIN la_oenb[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2300.870 -4.800 2301.430 1.000 ;
    END
  END la_oenb[98]
  PIN la_oenb[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2317.430 -4.800 2317.990 1.000 ;
    END
  END la_oenb[99]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 827.030 -4.800 827.590 1.000 ;
    END
  END la_oenb[9]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 8.970 10.640 12.070 3468.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 188.970 10.640 192.070 1260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 188.970 1696.540 192.070 1820.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 188.970 2256.540 192.070 2380.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 188.970 2816.540 192.070 2940.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 188.970 3376.540 192.070 3468.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 368.970 10.640 372.070 1260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 368.970 1696.540 372.070 1820.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 368.970 2256.540 372.070 2380.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 368.970 2816.540 372.070 2940.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 368.970 3376.540 372.070 3468.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 548.970 10.640 552.070 1260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 548.970 1696.540 552.070 1820.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 548.970 2256.540 552.070 2380.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 548.970 2816.540 552.070 2940.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 548.970 3376.540 552.070 3468.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 728.970 10.640 732.070 1260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 728.970 1696.540 732.070 1820.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 728.970 2256.540 732.070 2380.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 728.970 2816.540 732.070 2940.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 728.970 3376.540 732.070 3468.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 908.970 10.640 912.070 2940.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 908.970 3357.500 912.070 3468.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 1088.970 10.640 1092.070 2940.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1088.970 3357.500 1092.070 3468.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 1268.970 10.640 1272.070 2940.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1268.970 3357.500 1272.070 3468.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 1448.970 10.640 1452.070 3468.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 1628.970 10.640 1632.070 140.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1628.970 557.500 1632.070 2940.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1628.970 3357.500 1632.070 3468.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 1808.970 10.640 1812.070 140.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1808.970 557.500 1812.070 2940.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1808.970 3357.500 1812.070 3468.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 1988.970 10.640 1992.070 3468.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 2168.970 10.640 2172.070 140.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2168.970 576.540 2172.070 700.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2168.970 1136.540 2172.070 1260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2168.970 1696.540 2172.070 1820.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2168.970 2256.540 2172.070 2380.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2168.970 2816.540 2172.070 2940.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2168.970 3376.540 2172.070 3468.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 2348.970 10.640 2352.070 140.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2348.970 576.540 2352.070 700.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2348.970 1136.540 2352.070 1260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2348.970 1696.540 2352.070 1820.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2348.970 2256.540 2352.070 2380.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2348.970 2816.540 2352.070 2940.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2348.970 3376.540 2352.070 3468.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 2528.970 10.640 2532.070 140.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2528.970 576.540 2532.070 700.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2528.970 1136.540 2532.070 1260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2528.970 1696.540 2532.070 1820.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2528.970 2256.540 2532.070 2380.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2528.970 2816.540 2532.070 2940.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2528.970 3376.540 2532.070 3468.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 2708.970 10.640 2712.070 140.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2708.970 576.540 2712.070 700.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2708.970 1136.540 2712.070 1260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2708.970 1696.540 2712.070 1820.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2708.970 2256.540 2712.070 2380.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2708.970 2816.540 2712.070 2940.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2708.970 3376.540 2712.070 3468.240 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 14.330 2874.320 17.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 194.330 2874.320 197.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 374.330 2874.320 377.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 554.330 2874.320 557.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 734.330 2874.320 737.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 914.330 2874.320 917.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1094.330 2874.320 1097.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1274.330 2874.320 1277.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1454.330 2874.320 1457.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1634.330 2874.320 1637.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1814.330 2874.320 1817.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1994.330 2874.320 1997.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 2174.330 2874.320 2177.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 2354.330 2874.320 2357.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 2534.330 2874.320 2537.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 2714.330 2874.320 2717.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 2894.330 2874.320 2897.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 3074.330 2874.320 3077.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 3254.330 2874.320 3257.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 3434.330 2874.320 3437.430 ;
    END
    PORT
      LAYER met4 ;
        RECT 845.310 2934.640 848.410 3359.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 2831.590 138.480 2834.690 579.600 ;
    END
    PORT
      LAYER met4 ;
        RECT 2831.590 698.800 2834.690 1139.920 ;
    END
    PORT
      LAYER met4 ;
        RECT 2831.590 1259.120 2834.690 1700.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 2831.590 1819.440 2834.690 2260.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 2831.590 2379.760 2834.690 2820.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 2831.590 2934.640 2834.690 3381.200 ;
    END
    PORT
      LAYER met5 ;
        RECT 1988.970 635.950 2874.320 639.050 ;
    END
    PORT
      LAYER met5 ;
        RECT 1988.970 1196.950 2874.320 1200.050 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 98.970 10.640 102.070 1260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 98.970 1696.540 102.070 1820.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 98.970 2256.540 102.070 2380.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 98.970 2816.540 102.070 2940.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 98.970 3376.540 102.070 3468.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 278.970 10.640 282.070 1260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 278.970 1696.540 282.070 1820.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 278.970 2256.540 282.070 2380.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 278.970 2816.540 282.070 2940.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 278.970 3376.540 282.070 3468.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 458.970 10.640 462.070 1260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 458.970 1696.540 462.070 1820.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 458.970 2256.540 462.070 2380.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 458.970 2816.540 462.070 2940.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 458.970 3376.540 462.070 3468.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 638.970 10.640 642.070 1260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 638.970 1696.540 642.070 1820.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 638.970 2256.540 642.070 2380.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 638.970 2816.540 642.070 2940.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 638.970 3376.540 642.070 3468.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 818.970 10.640 822.070 3468.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 998.970 10.640 1002.070 2940.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 998.970 3357.500 1002.070 3468.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 1178.970 10.640 1182.070 2940.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1178.970 3357.500 1182.070 3468.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 1358.970 10.640 1362.070 2940.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1358.970 3357.500 1362.070 3468.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 1538.970 10.640 1542.070 140.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1538.970 557.500 1542.070 2940.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1538.970 3357.500 1542.070 3468.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 1718.970 10.640 1722.070 140.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1718.970 557.500 1722.070 2940.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1718.970 3357.500 1722.070 3468.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 1898.970 10.640 1902.070 140.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1898.970 557.500 1902.070 2940.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1898.970 3357.500 1902.070 3468.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 2078.970 10.640 2082.070 3468.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 2258.970 10.640 2262.070 140.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2258.970 576.540 2262.070 700.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2258.970 1136.540 2262.070 1260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2258.970 1696.540 2262.070 1820.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2258.970 2256.540 2262.070 2380.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2258.970 2816.540 2262.070 2940.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2258.970 3376.540 2262.070 3468.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 2438.970 10.640 2442.070 140.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2438.970 576.540 2442.070 700.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2438.970 1136.540 2442.070 1260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2438.970 1696.540 2442.070 1820.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2438.970 2256.540 2442.070 2380.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2438.970 2816.540 2442.070 2940.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2438.970 3376.540 2442.070 3468.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 2618.970 10.640 2622.070 140.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2618.970 576.540 2622.070 700.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2618.970 1136.540 2622.070 1260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2618.970 1696.540 2622.070 1820.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2618.970 2256.540 2622.070 2380.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2618.970 2816.540 2622.070 2940.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2618.970 3376.540 2622.070 3468.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 2798.970 10.640 2802.070 3468.240 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 104.330 2874.320 107.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 284.330 2874.320 287.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 464.330 2874.320 467.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 644.330 2874.320 647.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 824.330 2874.320 827.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1004.330 2874.320 1007.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1184.330 2874.320 1187.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1364.330 2874.320 1367.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1544.330 2874.320 1547.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1724.330 2874.320 1727.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 1904.330 2874.320 1907.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 2084.330 2874.320 2087.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 2264.330 2874.320 2267.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 2444.330 2874.320 2447.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 2624.330 2874.320 2627.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 2804.330 2874.320 2807.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 2984.330 2874.320 2987.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 3164.330 2874.320 3167.430 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 3344.330 2874.320 3347.430 ;
    END
    PORT
      LAYER met4 ;
        RECT 45.830 1256.400 48.930 1697.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 45.830 1816.720 48.930 2257.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 1437.790 2937.360 1440.890 3362.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 45.830 2377.040 48.930 2818.160 ;
    END
    PORT
      LAYER met5 ;
        RECT 818.970 3410.350 2082.070 3413.450 ;
    END
    PORT
      LAYER met4 ;
        RECT 45.830 2937.360 48.930 3378.480 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 3420.550 822.070 3423.650 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 2876.550 822.070 2879.650 ;
    END
    PORT
      LAYER met5 ;
        RECT 2078.970 2876.550 2802.070 2879.650 ;
    END
    PORT
      LAYER met5 ;
        RECT 2078.970 3420.550 2802.070 3423.650 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.830 -4.800 82.390 1.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.350 -4.800 87.910 1.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.870 -4.800 93.430 1.000 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 114.950 -4.800 115.510 1.000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 302.630 -4.800 303.190 1.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 319.190 -4.800 319.750 1.000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 335.750 -4.800 336.310 1.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 352.310 -4.800 352.870 1.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 368.870 -4.800 369.430 1.000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 385.430 -4.800 385.990 1.000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 401.990 -4.800 402.550 1.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 418.550 -4.800 419.110 1.000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 435.110 -4.800 435.670 1.000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 451.670 -4.800 452.230 1.000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 137.030 -4.800 137.590 1.000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 468.230 -4.800 468.790 1.000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 484.790 -4.800 485.350 1.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 501.350 -4.800 501.910 1.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 517.910 -4.800 518.470 1.000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 534.470 -4.800 535.030 1.000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 551.030 -4.800 551.590 1.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 567.590 -4.800 568.150 1.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 584.150 -4.800 584.710 1.000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 600.710 -4.800 601.270 1.000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 617.270 -4.800 617.830 1.000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 159.110 -4.800 159.670 1.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 633.830 -4.800 634.390 1.000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 650.390 -4.800 650.950 1.000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 181.190 -4.800 181.750 1.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 203.270 -4.800 203.830 1.000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.830 -4.800 220.390 1.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.390 -4.800 236.950 1.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 252.950 -4.800 253.510 1.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 269.510 -4.800 270.070 1.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.070 -4.800 286.630 1.000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.390 -4.800 98.950 1.000 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.470 -4.800 121.030 1.000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 308.150 -4.800 308.710 1.000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 324.710 -4.800 325.270 1.000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 341.270 -4.800 341.830 1.000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.830 -4.800 358.390 1.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 374.390 -4.800 374.950 1.000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 390.950 -4.800 391.510 1.000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 407.510 -4.800 408.070 1.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 424.070 -4.800 424.630 1.000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 440.630 -4.800 441.190 1.000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 457.190 -4.800 457.750 1.000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 142.550 -4.800 143.110 1.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 473.750 -4.800 474.310 1.000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 490.310 -4.800 490.870 1.000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 506.870 -4.800 507.430 1.000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 523.430 -4.800 523.990 1.000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 539.990 -4.800 540.550 1.000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 556.550 -4.800 557.110 1.000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 573.110 -4.800 573.670 1.000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 589.670 -4.800 590.230 1.000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 606.230 -4.800 606.790 1.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 622.790 -4.800 623.350 1.000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.630 -4.800 165.190 1.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 639.350 -4.800 639.910 1.000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 655.910 -4.800 656.470 1.000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.710 -4.800 187.270 1.000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.790 -4.800 209.350 1.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.350 -4.800 225.910 1.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.910 -4.800 242.470 1.000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 258.470 -4.800 259.030 1.000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 275.030 -4.800 275.590 1.000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 291.590 -4.800 292.150 1.000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.990 -4.800 126.550 1.000 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 313.670 -4.800 314.230 1.000 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 330.230 -4.800 330.790 1.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 346.790 -4.800 347.350 1.000 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.350 -4.800 363.910 1.000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 379.910 -4.800 380.470 1.000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 396.470 -4.800 397.030 1.000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 413.030 -4.800 413.590 1.000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 429.590 -4.800 430.150 1.000 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 446.150 -4.800 446.710 1.000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 462.710 -4.800 463.270 1.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.070 -4.800 148.630 1.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 479.270 -4.800 479.830 1.000 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 495.830 -4.800 496.390 1.000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 512.390 -4.800 512.950 1.000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 528.950 -4.800 529.510 1.000 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 545.510 -4.800 546.070 1.000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 562.070 -4.800 562.630 1.000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 578.630 -4.800 579.190 1.000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 595.190 -4.800 595.750 1.000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 611.750 -4.800 612.310 1.000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 628.310 -4.800 628.870 1.000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.150 -4.800 170.710 1.000 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 644.870 -4.800 645.430 1.000 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 661.430 -4.800 661.990 1.000 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 192.230 -4.800 192.790 1.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 214.310 -4.800 214.870 1.000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 230.870 -4.800 231.430 1.000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 247.430 -4.800 247.990 1.000 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 263.990 -4.800 264.550 1.000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.550 -4.800 281.110 1.000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 297.110 -4.800 297.670 1.000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.510 -4.800 132.070 1.000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 153.590 -4.800 154.150 1.000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 175.670 -4.800 176.230 1.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 197.750 -4.800 198.310 1.000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.910 -4.800 104.470 1.000 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.430 -4.800 109.990 1.000 ;
    END
  END wbs_we_i
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 2874.080 3468.085 ;
      LAYER met1 ;
        RECT 3.750 6.840 2874.080 3468.240 ;
      LAYER met2 ;
        RECT 3.770 3478.720 58.090 3479.290 ;
        RECT 59.210 3478.720 164.350 3479.290 ;
        RECT 165.470 3478.720 270.610 3479.290 ;
        RECT 271.730 3478.720 376.870 3479.290 ;
        RECT 377.990 3478.720 483.130 3479.290 ;
        RECT 484.250 3478.720 589.390 3479.290 ;
        RECT 590.510 3478.720 695.650 3479.290 ;
        RECT 696.770 3478.720 801.910 3479.290 ;
        RECT 803.030 3478.720 908.170 3479.290 ;
        RECT 909.290 3478.720 1014.430 3479.290 ;
        RECT 1015.550 3478.720 1120.690 3479.290 ;
        RECT 1121.810 3478.720 1226.950 3479.290 ;
        RECT 1228.070 3478.720 1333.210 3479.290 ;
        RECT 1334.330 3478.720 1439.470 3479.290 ;
        RECT 1440.590 3478.720 1545.730 3479.290 ;
        RECT 1546.850 3478.720 1651.990 3479.290 ;
        RECT 1653.110 3478.720 1758.250 3479.290 ;
        RECT 1759.370 3478.720 1864.510 3479.290 ;
        RECT 1865.630 3478.720 1970.770 3479.290 ;
        RECT 1971.890 3478.720 2077.030 3479.290 ;
        RECT 2078.150 3478.720 2183.290 3479.290 ;
        RECT 2184.410 3478.720 2289.550 3479.290 ;
        RECT 2290.670 3478.720 2395.810 3479.290 ;
        RECT 2396.930 3478.720 2502.070 3479.290 ;
        RECT 2503.190 3478.720 2608.330 3479.290 ;
        RECT 2609.450 3478.720 2714.590 3479.290 ;
        RECT 2715.710 3478.720 2820.850 3479.290 ;
        RECT 2821.970 3478.720 2870.770 3479.290 ;
        RECT 3.770 1.280 2870.770 3478.720 ;
        RECT 3.770 0.270 81.550 1.280 ;
        RECT 82.670 0.270 87.070 1.280 ;
        RECT 88.190 0.270 92.590 1.280 ;
        RECT 93.710 0.270 98.110 1.280 ;
        RECT 99.230 0.270 103.630 1.280 ;
        RECT 104.750 0.270 109.150 1.280 ;
        RECT 110.270 0.270 114.670 1.280 ;
        RECT 115.790 0.270 120.190 1.280 ;
        RECT 121.310 0.270 125.710 1.280 ;
        RECT 126.830 0.270 131.230 1.280 ;
        RECT 132.350 0.270 136.750 1.280 ;
        RECT 137.870 0.270 142.270 1.280 ;
        RECT 143.390 0.270 147.790 1.280 ;
        RECT 148.910 0.270 153.310 1.280 ;
        RECT 154.430 0.270 158.830 1.280 ;
        RECT 159.950 0.270 164.350 1.280 ;
        RECT 165.470 0.270 169.870 1.280 ;
        RECT 170.990 0.270 175.390 1.280 ;
        RECT 176.510 0.270 180.910 1.280 ;
        RECT 182.030 0.270 186.430 1.280 ;
        RECT 187.550 0.270 191.950 1.280 ;
        RECT 193.070 0.270 197.470 1.280 ;
        RECT 198.590 0.270 202.990 1.280 ;
        RECT 204.110 0.270 208.510 1.280 ;
        RECT 209.630 0.270 214.030 1.280 ;
        RECT 215.150 0.270 219.550 1.280 ;
        RECT 220.670 0.270 225.070 1.280 ;
        RECT 226.190 0.270 230.590 1.280 ;
        RECT 231.710 0.270 236.110 1.280 ;
        RECT 237.230 0.270 241.630 1.280 ;
        RECT 242.750 0.270 247.150 1.280 ;
        RECT 248.270 0.270 252.670 1.280 ;
        RECT 253.790 0.270 258.190 1.280 ;
        RECT 259.310 0.270 263.710 1.280 ;
        RECT 264.830 0.270 269.230 1.280 ;
        RECT 270.350 0.270 274.750 1.280 ;
        RECT 275.870 0.270 280.270 1.280 ;
        RECT 281.390 0.270 285.790 1.280 ;
        RECT 286.910 0.270 291.310 1.280 ;
        RECT 292.430 0.270 296.830 1.280 ;
        RECT 297.950 0.270 302.350 1.280 ;
        RECT 303.470 0.270 307.870 1.280 ;
        RECT 308.990 0.270 313.390 1.280 ;
        RECT 314.510 0.270 318.910 1.280 ;
        RECT 320.030 0.270 324.430 1.280 ;
        RECT 325.550 0.270 329.950 1.280 ;
        RECT 331.070 0.270 335.470 1.280 ;
        RECT 336.590 0.270 340.990 1.280 ;
        RECT 342.110 0.270 346.510 1.280 ;
        RECT 347.630 0.270 352.030 1.280 ;
        RECT 353.150 0.270 357.550 1.280 ;
        RECT 358.670 0.270 363.070 1.280 ;
        RECT 364.190 0.270 368.590 1.280 ;
        RECT 369.710 0.270 374.110 1.280 ;
        RECT 375.230 0.270 379.630 1.280 ;
        RECT 380.750 0.270 385.150 1.280 ;
        RECT 386.270 0.270 390.670 1.280 ;
        RECT 391.790 0.270 396.190 1.280 ;
        RECT 397.310 0.270 401.710 1.280 ;
        RECT 402.830 0.270 407.230 1.280 ;
        RECT 408.350 0.270 412.750 1.280 ;
        RECT 413.870 0.270 418.270 1.280 ;
        RECT 419.390 0.270 423.790 1.280 ;
        RECT 424.910 0.270 429.310 1.280 ;
        RECT 430.430 0.270 434.830 1.280 ;
        RECT 435.950 0.270 440.350 1.280 ;
        RECT 441.470 0.270 445.870 1.280 ;
        RECT 446.990 0.270 451.390 1.280 ;
        RECT 452.510 0.270 456.910 1.280 ;
        RECT 458.030 0.270 462.430 1.280 ;
        RECT 463.550 0.270 467.950 1.280 ;
        RECT 469.070 0.270 473.470 1.280 ;
        RECT 474.590 0.270 478.990 1.280 ;
        RECT 480.110 0.270 484.510 1.280 ;
        RECT 485.630 0.270 490.030 1.280 ;
        RECT 491.150 0.270 495.550 1.280 ;
        RECT 496.670 0.270 501.070 1.280 ;
        RECT 502.190 0.270 506.590 1.280 ;
        RECT 507.710 0.270 512.110 1.280 ;
        RECT 513.230 0.270 517.630 1.280 ;
        RECT 518.750 0.270 523.150 1.280 ;
        RECT 524.270 0.270 528.670 1.280 ;
        RECT 529.790 0.270 534.190 1.280 ;
        RECT 535.310 0.270 539.710 1.280 ;
        RECT 540.830 0.270 545.230 1.280 ;
        RECT 546.350 0.270 550.750 1.280 ;
        RECT 551.870 0.270 556.270 1.280 ;
        RECT 557.390 0.270 561.790 1.280 ;
        RECT 562.910 0.270 567.310 1.280 ;
        RECT 568.430 0.270 572.830 1.280 ;
        RECT 573.950 0.270 578.350 1.280 ;
        RECT 579.470 0.270 583.870 1.280 ;
        RECT 584.990 0.270 589.390 1.280 ;
        RECT 590.510 0.270 594.910 1.280 ;
        RECT 596.030 0.270 600.430 1.280 ;
        RECT 601.550 0.270 605.950 1.280 ;
        RECT 607.070 0.270 611.470 1.280 ;
        RECT 612.590 0.270 616.990 1.280 ;
        RECT 618.110 0.270 622.510 1.280 ;
        RECT 623.630 0.270 628.030 1.280 ;
        RECT 629.150 0.270 633.550 1.280 ;
        RECT 634.670 0.270 639.070 1.280 ;
        RECT 640.190 0.270 644.590 1.280 ;
        RECT 645.710 0.270 650.110 1.280 ;
        RECT 651.230 0.270 655.630 1.280 ;
        RECT 656.750 0.270 661.150 1.280 ;
        RECT 662.270 0.270 666.670 1.280 ;
        RECT 667.790 0.270 672.190 1.280 ;
        RECT 673.310 0.270 677.710 1.280 ;
        RECT 678.830 0.270 683.230 1.280 ;
        RECT 684.350 0.270 688.750 1.280 ;
        RECT 689.870 0.270 694.270 1.280 ;
        RECT 695.390 0.270 699.790 1.280 ;
        RECT 700.910 0.270 705.310 1.280 ;
        RECT 706.430 0.270 710.830 1.280 ;
        RECT 711.950 0.270 716.350 1.280 ;
        RECT 717.470 0.270 721.870 1.280 ;
        RECT 722.990 0.270 727.390 1.280 ;
        RECT 728.510 0.270 732.910 1.280 ;
        RECT 734.030 0.270 738.430 1.280 ;
        RECT 739.550 0.270 743.950 1.280 ;
        RECT 745.070 0.270 749.470 1.280 ;
        RECT 750.590 0.270 754.990 1.280 ;
        RECT 756.110 0.270 760.510 1.280 ;
        RECT 761.630 0.270 766.030 1.280 ;
        RECT 767.150 0.270 771.550 1.280 ;
        RECT 772.670 0.270 777.070 1.280 ;
        RECT 778.190 0.270 782.590 1.280 ;
        RECT 783.710 0.270 788.110 1.280 ;
        RECT 789.230 0.270 793.630 1.280 ;
        RECT 794.750 0.270 799.150 1.280 ;
        RECT 800.270 0.270 804.670 1.280 ;
        RECT 805.790 0.270 810.190 1.280 ;
        RECT 811.310 0.270 815.710 1.280 ;
        RECT 816.830 0.270 821.230 1.280 ;
        RECT 822.350 0.270 826.750 1.280 ;
        RECT 827.870 0.270 832.270 1.280 ;
        RECT 833.390 0.270 837.790 1.280 ;
        RECT 838.910 0.270 843.310 1.280 ;
        RECT 844.430 0.270 848.830 1.280 ;
        RECT 849.950 0.270 854.350 1.280 ;
        RECT 855.470 0.270 859.870 1.280 ;
        RECT 860.990 0.270 865.390 1.280 ;
        RECT 866.510 0.270 870.910 1.280 ;
        RECT 872.030 0.270 876.430 1.280 ;
        RECT 877.550 0.270 881.950 1.280 ;
        RECT 883.070 0.270 887.470 1.280 ;
        RECT 888.590 0.270 892.990 1.280 ;
        RECT 894.110 0.270 898.510 1.280 ;
        RECT 899.630 0.270 904.030 1.280 ;
        RECT 905.150 0.270 909.550 1.280 ;
        RECT 910.670 0.270 915.070 1.280 ;
        RECT 916.190 0.270 920.590 1.280 ;
        RECT 921.710 0.270 926.110 1.280 ;
        RECT 927.230 0.270 931.630 1.280 ;
        RECT 932.750 0.270 937.150 1.280 ;
        RECT 938.270 0.270 942.670 1.280 ;
        RECT 943.790 0.270 948.190 1.280 ;
        RECT 949.310 0.270 953.710 1.280 ;
        RECT 954.830 0.270 959.230 1.280 ;
        RECT 960.350 0.270 964.750 1.280 ;
        RECT 965.870 0.270 970.270 1.280 ;
        RECT 971.390 0.270 975.790 1.280 ;
        RECT 976.910 0.270 981.310 1.280 ;
        RECT 982.430 0.270 986.830 1.280 ;
        RECT 987.950 0.270 992.350 1.280 ;
        RECT 993.470 0.270 997.870 1.280 ;
        RECT 998.990 0.270 1003.390 1.280 ;
        RECT 1004.510 0.270 1008.910 1.280 ;
        RECT 1010.030 0.270 1014.430 1.280 ;
        RECT 1015.550 0.270 1019.950 1.280 ;
        RECT 1021.070 0.270 1025.470 1.280 ;
        RECT 1026.590 0.270 1030.990 1.280 ;
        RECT 1032.110 0.270 1036.510 1.280 ;
        RECT 1037.630 0.270 1042.030 1.280 ;
        RECT 1043.150 0.270 1047.550 1.280 ;
        RECT 1048.670 0.270 1053.070 1.280 ;
        RECT 1054.190 0.270 1058.590 1.280 ;
        RECT 1059.710 0.270 1064.110 1.280 ;
        RECT 1065.230 0.270 1069.630 1.280 ;
        RECT 1070.750 0.270 1075.150 1.280 ;
        RECT 1076.270 0.270 1080.670 1.280 ;
        RECT 1081.790 0.270 1086.190 1.280 ;
        RECT 1087.310 0.270 1091.710 1.280 ;
        RECT 1092.830 0.270 1097.230 1.280 ;
        RECT 1098.350 0.270 1102.750 1.280 ;
        RECT 1103.870 0.270 1108.270 1.280 ;
        RECT 1109.390 0.270 1113.790 1.280 ;
        RECT 1114.910 0.270 1119.310 1.280 ;
        RECT 1120.430 0.270 1124.830 1.280 ;
        RECT 1125.950 0.270 1130.350 1.280 ;
        RECT 1131.470 0.270 1135.870 1.280 ;
        RECT 1136.990 0.270 1141.390 1.280 ;
        RECT 1142.510 0.270 1146.910 1.280 ;
        RECT 1148.030 0.270 1152.430 1.280 ;
        RECT 1153.550 0.270 1157.950 1.280 ;
        RECT 1159.070 0.270 1163.470 1.280 ;
        RECT 1164.590 0.270 1168.990 1.280 ;
        RECT 1170.110 0.270 1174.510 1.280 ;
        RECT 1175.630 0.270 1180.030 1.280 ;
        RECT 1181.150 0.270 1185.550 1.280 ;
        RECT 1186.670 0.270 1191.070 1.280 ;
        RECT 1192.190 0.270 1196.590 1.280 ;
        RECT 1197.710 0.270 1202.110 1.280 ;
        RECT 1203.230 0.270 1207.630 1.280 ;
        RECT 1208.750 0.270 1213.150 1.280 ;
        RECT 1214.270 0.270 1218.670 1.280 ;
        RECT 1219.790 0.270 1224.190 1.280 ;
        RECT 1225.310 0.270 1229.710 1.280 ;
        RECT 1230.830 0.270 1235.230 1.280 ;
        RECT 1236.350 0.270 1240.750 1.280 ;
        RECT 1241.870 0.270 1246.270 1.280 ;
        RECT 1247.390 0.270 1251.790 1.280 ;
        RECT 1252.910 0.270 1257.310 1.280 ;
        RECT 1258.430 0.270 1262.830 1.280 ;
        RECT 1263.950 0.270 1268.350 1.280 ;
        RECT 1269.470 0.270 1273.870 1.280 ;
        RECT 1274.990 0.270 1279.390 1.280 ;
        RECT 1280.510 0.270 1284.910 1.280 ;
        RECT 1286.030 0.270 1290.430 1.280 ;
        RECT 1291.550 0.270 1295.950 1.280 ;
        RECT 1297.070 0.270 1301.470 1.280 ;
        RECT 1302.590 0.270 1306.990 1.280 ;
        RECT 1308.110 0.270 1312.510 1.280 ;
        RECT 1313.630 0.270 1318.030 1.280 ;
        RECT 1319.150 0.270 1323.550 1.280 ;
        RECT 1324.670 0.270 1329.070 1.280 ;
        RECT 1330.190 0.270 1334.590 1.280 ;
        RECT 1335.710 0.270 1340.110 1.280 ;
        RECT 1341.230 0.270 1345.630 1.280 ;
        RECT 1346.750 0.270 1351.150 1.280 ;
        RECT 1352.270 0.270 1356.670 1.280 ;
        RECT 1357.790 0.270 1362.190 1.280 ;
        RECT 1363.310 0.270 1367.710 1.280 ;
        RECT 1368.830 0.270 1373.230 1.280 ;
        RECT 1374.350 0.270 1378.750 1.280 ;
        RECT 1379.870 0.270 1384.270 1.280 ;
        RECT 1385.390 0.270 1389.790 1.280 ;
        RECT 1390.910 0.270 1395.310 1.280 ;
        RECT 1396.430 0.270 1400.830 1.280 ;
        RECT 1401.950 0.270 1406.350 1.280 ;
        RECT 1407.470 0.270 1411.870 1.280 ;
        RECT 1412.990 0.270 1417.390 1.280 ;
        RECT 1418.510 0.270 1422.910 1.280 ;
        RECT 1424.030 0.270 1428.430 1.280 ;
        RECT 1429.550 0.270 1433.950 1.280 ;
        RECT 1435.070 0.270 1439.470 1.280 ;
        RECT 1440.590 0.270 1444.990 1.280 ;
        RECT 1446.110 0.270 1450.510 1.280 ;
        RECT 1451.630 0.270 1456.030 1.280 ;
        RECT 1457.150 0.270 1461.550 1.280 ;
        RECT 1462.670 0.270 1467.070 1.280 ;
        RECT 1468.190 0.270 1472.590 1.280 ;
        RECT 1473.710 0.270 1478.110 1.280 ;
        RECT 1479.230 0.270 1483.630 1.280 ;
        RECT 1484.750 0.270 1489.150 1.280 ;
        RECT 1490.270 0.270 1494.670 1.280 ;
        RECT 1495.790 0.270 1500.190 1.280 ;
        RECT 1501.310 0.270 1505.710 1.280 ;
        RECT 1506.830 0.270 1511.230 1.280 ;
        RECT 1512.350 0.270 1516.750 1.280 ;
        RECT 1517.870 0.270 1522.270 1.280 ;
        RECT 1523.390 0.270 1527.790 1.280 ;
        RECT 1528.910 0.270 1533.310 1.280 ;
        RECT 1534.430 0.270 1538.830 1.280 ;
        RECT 1539.950 0.270 1544.350 1.280 ;
        RECT 1545.470 0.270 1549.870 1.280 ;
        RECT 1550.990 0.270 1555.390 1.280 ;
        RECT 1556.510 0.270 1560.910 1.280 ;
        RECT 1562.030 0.270 1566.430 1.280 ;
        RECT 1567.550 0.270 1571.950 1.280 ;
        RECT 1573.070 0.270 1577.470 1.280 ;
        RECT 1578.590 0.270 1582.990 1.280 ;
        RECT 1584.110 0.270 1588.510 1.280 ;
        RECT 1589.630 0.270 1594.030 1.280 ;
        RECT 1595.150 0.270 1599.550 1.280 ;
        RECT 1600.670 0.270 1605.070 1.280 ;
        RECT 1606.190 0.270 1610.590 1.280 ;
        RECT 1611.710 0.270 1616.110 1.280 ;
        RECT 1617.230 0.270 1621.630 1.280 ;
        RECT 1622.750 0.270 1627.150 1.280 ;
        RECT 1628.270 0.270 1632.670 1.280 ;
        RECT 1633.790 0.270 1638.190 1.280 ;
        RECT 1639.310 0.270 1643.710 1.280 ;
        RECT 1644.830 0.270 1649.230 1.280 ;
        RECT 1650.350 0.270 1654.750 1.280 ;
        RECT 1655.870 0.270 1660.270 1.280 ;
        RECT 1661.390 0.270 1665.790 1.280 ;
        RECT 1666.910 0.270 1671.310 1.280 ;
        RECT 1672.430 0.270 1676.830 1.280 ;
        RECT 1677.950 0.270 1682.350 1.280 ;
        RECT 1683.470 0.270 1687.870 1.280 ;
        RECT 1688.990 0.270 1693.390 1.280 ;
        RECT 1694.510 0.270 1698.910 1.280 ;
        RECT 1700.030 0.270 1704.430 1.280 ;
        RECT 1705.550 0.270 1709.950 1.280 ;
        RECT 1711.070 0.270 1715.470 1.280 ;
        RECT 1716.590 0.270 1720.990 1.280 ;
        RECT 1722.110 0.270 1726.510 1.280 ;
        RECT 1727.630 0.270 1732.030 1.280 ;
        RECT 1733.150 0.270 1737.550 1.280 ;
        RECT 1738.670 0.270 1743.070 1.280 ;
        RECT 1744.190 0.270 1748.590 1.280 ;
        RECT 1749.710 0.270 1754.110 1.280 ;
        RECT 1755.230 0.270 1759.630 1.280 ;
        RECT 1760.750 0.270 1765.150 1.280 ;
        RECT 1766.270 0.270 1770.670 1.280 ;
        RECT 1771.790 0.270 1776.190 1.280 ;
        RECT 1777.310 0.270 1781.710 1.280 ;
        RECT 1782.830 0.270 1787.230 1.280 ;
        RECT 1788.350 0.270 1792.750 1.280 ;
        RECT 1793.870 0.270 1798.270 1.280 ;
        RECT 1799.390 0.270 1803.790 1.280 ;
        RECT 1804.910 0.270 1809.310 1.280 ;
        RECT 1810.430 0.270 1814.830 1.280 ;
        RECT 1815.950 0.270 1820.350 1.280 ;
        RECT 1821.470 0.270 1825.870 1.280 ;
        RECT 1826.990 0.270 1831.390 1.280 ;
        RECT 1832.510 0.270 1836.910 1.280 ;
        RECT 1838.030 0.270 1842.430 1.280 ;
        RECT 1843.550 0.270 1847.950 1.280 ;
        RECT 1849.070 0.270 1853.470 1.280 ;
        RECT 1854.590 0.270 1858.990 1.280 ;
        RECT 1860.110 0.270 1864.510 1.280 ;
        RECT 1865.630 0.270 1870.030 1.280 ;
        RECT 1871.150 0.270 1875.550 1.280 ;
        RECT 1876.670 0.270 1881.070 1.280 ;
        RECT 1882.190 0.270 1886.590 1.280 ;
        RECT 1887.710 0.270 1892.110 1.280 ;
        RECT 1893.230 0.270 1897.630 1.280 ;
        RECT 1898.750 0.270 1903.150 1.280 ;
        RECT 1904.270 0.270 1908.670 1.280 ;
        RECT 1909.790 0.270 1914.190 1.280 ;
        RECT 1915.310 0.270 1919.710 1.280 ;
        RECT 1920.830 0.270 1925.230 1.280 ;
        RECT 1926.350 0.270 1930.750 1.280 ;
        RECT 1931.870 0.270 1936.270 1.280 ;
        RECT 1937.390 0.270 1941.790 1.280 ;
        RECT 1942.910 0.270 1947.310 1.280 ;
        RECT 1948.430 0.270 1952.830 1.280 ;
        RECT 1953.950 0.270 1958.350 1.280 ;
        RECT 1959.470 0.270 1963.870 1.280 ;
        RECT 1964.990 0.270 1969.390 1.280 ;
        RECT 1970.510 0.270 1974.910 1.280 ;
        RECT 1976.030 0.270 1980.430 1.280 ;
        RECT 1981.550 0.270 1985.950 1.280 ;
        RECT 1987.070 0.270 1991.470 1.280 ;
        RECT 1992.590 0.270 1996.990 1.280 ;
        RECT 1998.110 0.270 2002.510 1.280 ;
        RECT 2003.630 0.270 2008.030 1.280 ;
        RECT 2009.150 0.270 2013.550 1.280 ;
        RECT 2014.670 0.270 2019.070 1.280 ;
        RECT 2020.190 0.270 2024.590 1.280 ;
        RECT 2025.710 0.270 2030.110 1.280 ;
        RECT 2031.230 0.270 2035.630 1.280 ;
        RECT 2036.750 0.270 2041.150 1.280 ;
        RECT 2042.270 0.270 2046.670 1.280 ;
        RECT 2047.790 0.270 2052.190 1.280 ;
        RECT 2053.310 0.270 2057.710 1.280 ;
        RECT 2058.830 0.270 2063.230 1.280 ;
        RECT 2064.350 0.270 2068.750 1.280 ;
        RECT 2069.870 0.270 2074.270 1.280 ;
        RECT 2075.390 0.270 2079.790 1.280 ;
        RECT 2080.910 0.270 2085.310 1.280 ;
        RECT 2086.430 0.270 2090.830 1.280 ;
        RECT 2091.950 0.270 2096.350 1.280 ;
        RECT 2097.470 0.270 2101.870 1.280 ;
        RECT 2102.990 0.270 2107.390 1.280 ;
        RECT 2108.510 0.270 2112.910 1.280 ;
        RECT 2114.030 0.270 2118.430 1.280 ;
        RECT 2119.550 0.270 2123.950 1.280 ;
        RECT 2125.070 0.270 2129.470 1.280 ;
        RECT 2130.590 0.270 2134.990 1.280 ;
        RECT 2136.110 0.270 2140.510 1.280 ;
        RECT 2141.630 0.270 2146.030 1.280 ;
        RECT 2147.150 0.270 2151.550 1.280 ;
        RECT 2152.670 0.270 2157.070 1.280 ;
        RECT 2158.190 0.270 2162.590 1.280 ;
        RECT 2163.710 0.270 2168.110 1.280 ;
        RECT 2169.230 0.270 2173.630 1.280 ;
        RECT 2174.750 0.270 2179.150 1.280 ;
        RECT 2180.270 0.270 2184.670 1.280 ;
        RECT 2185.790 0.270 2190.190 1.280 ;
        RECT 2191.310 0.270 2195.710 1.280 ;
        RECT 2196.830 0.270 2201.230 1.280 ;
        RECT 2202.350 0.270 2206.750 1.280 ;
        RECT 2207.870 0.270 2212.270 1.280 ;
        RECT 2213.390 0.270 2217.790 1.280 ;
        RECT 2218.910 0.270 2223.310 1.280 ;
        RECT 2224.430 0.270 2228.830 1.280 ;
        RECT 2229.950 0.270 2234.350 1.280 ;
        RECT 2235.470 0.270 2239.870 1.280 ;
        RECT 2240.990 0.270 2245.390 1.280 ;
        RECT 2246.510 0.270 2250.910 1.280 ;
        RECT 2252.030 0.270 2256.430 1.280 ;
        RECT 2257.550 0.270 2261.950 1.280 ;
        RECT 2263.070 0.270 2267.470 1.280 ;
        RECT 2268.590 0.270 2272.990 1.280 ;
        RECT 2274.110 0.270 2278.510 1.280 ;
        RECT 2279.630 0.270 2284.030 1.280 ;
        RECT 2285.150 0.270 2289.550 1.280 ;
        RECT 2290.670 0.270 2295.070 1.280 ;
        RECT 2296.190 0.270 2300.590 1.280 ;
        RECT 2301.710 0.270 2306.110 1.280 ;
        RECT 2307.230 0.270 2311.630 1.280 ;
        RECT 2312.750 0.270 2317.150 1.280 ;
        RECT 2318.270 0.270 2322.670 1.280 ;
        RECT 2323.790 0.270 2328.190 1.280 ;
        RECT 2329.310 0.270 2333.710 1.280 ;
        RECT 2334.830 0.270 2339.230 1.280 ;
        RECT 2340.350 0.270 2344.750 1.280 ;
        RECT 2345.870 0.270 2350.270 1.280 ;
        RECT 2351.390 0.270 2355.790 1.280 ;
        RECT 2356.910 0.270 2361.310 1.280 ;
        RECT 2362.430 0.270 2366.830 1.280 ;
        RECT 2367.950 0.270 2372.350 1.280 ;
        RECT 2373.470 0.270 2377.870 1.280 ;
        RECT 2378.990 0.270 2383.390 1.280 ;
        RECT 2384.510 0.270 2388.910 1.280 ;
        RECT 2390.030 0.270 2394.430 1.280 ;
        RECT 2395.550 0.270 2399.950 1.280 ;
        RECT 2401.070 0.270 2405.470 1.280 ;
        RECT 2406.590 0.270 2410.990 1.280 ;
        RECT 2412.110 0.270 2416.510 1.280 ;
        RECT 2417.630 0.270 2422.030 1.280 ;
        RECT 2423.150 0.270 2427.550 1.280 ;
        RECT 2428.670 0.270 2433.070 1.280 ;
        RECT 2434.190 0.270 2438.590 1.280 ;
        RECT 2439.710 0.270 2444.110 1.280 ;
        RECT 2445.230 0.270 2449.630 1.280 ;
        RECT 2450.750 0.270 2455.150 1.280 ;
        RECT 2456.270 0.270 2460.670 1.280 ;
        RECT 2461.790 0.270 2466.190 1.280 ;
        RECT 2467.310 0.270 2471.710 1.280 ;
        RECT 2472.830 0.270 2477.230 1.280 ;
        RECT 2478.350 0.270 2482.750 1.280 ;
        RECT 2483.870 0.270 2488.270 1.280 ;
        RECT 2489.390 0.270 2493.790 1.280 ;
        RECT 2494.910 0.270 2499.310 1.280 ;
        RECT 2500.430 0.270 2504.830 1.280 ;
        RECT 2505.950 0.270 2510.350 1.280 ;
        RECT 2511.470 0.270 2515.870 1.280 ;
        RECT 2516.990 0.270 2521.390 1.280 ;
        RECT 2522.510 0.270 2526.910 1.280 ;
        RECT 2528.030 0.270 2532.430 1.280 ;
        RECT 2533.550 0.270 2537.950 1.280 ;
        RECT 2539.070 0.270 2543.470 1.280 ;
        RECT 2544.590 0.270 2548.990 1.280 ;
        RECT 2550.110 0.270 2554.510 1.280 ;
        RECT 2555.630 0.270 2560.030 1.280 ;
        RECT 2561.150 0.270 2565.550 1.280 ;
        RECT 2566.670 0.270 2571.070 1.280 ;
        RECT 2572.190 0.270 2576.590 1.280 ;
        RECT 2577.710 0.270 2582.110 1.280 ;
        RECT 2583.230 0.270 2587.630 1.280 ;
        RECT 2588.750 0.270 2593.150 1.280 ;
        RECT 2594.270 0.270 2598.670 1.280 ;
        RECT 2599.790 0.270 2604.190 1.280 ;
        RECT 2605.310 0.270 2609.710 1.280 ;
        RECT 2610.830 0.270 2615.230 1.280 ;
        RECT 2616.350 0.270 2620.750 1.280 ;
        RECT 2621.870 0.270 2626.270 1.280 ;
        RECT 2627.390 0.270 2631.790 1.280 ;
        RECT 2632.910 0.270 2637.310 1.280 ;
        RECT 2638.430 0.270 2642.830 1.280 ;
        RECT 2643.950 0.270 2648.350 1.280 ;
        RECT 2649.470 0.270 2653.870 1.280 ;
        RECT 2654.990 0.270 2659.390 1.280 ;
        RECT 2660.510 0.270 2664.910 1.280 ;
        RECT 2666.030 0.270 2670.430 1.280 ;
        RECT 2671.550 0.270 2675.950 1.280 ;
        RECT 2677.070 0.270 2681.470 1.280 ;
        RECT 2682.590 0.270 2686.990 1.280 ;
        RECT 2688.110 0.270 2692.510 1.280 ;
        RECT 2693.630 0.270 2698.030 1.280 ;
        RECT 2699.150 0.270 2703.550 1.280 ;
        RECT 2704.670 0.270 2709.070 1.280 ;
        RECT 2710.190 0.270 2714.590 1.280 ;
        RECT 2715.710 0.270 2720.110 1.280 ;
        RECT 2721.230 0.270 2725.630 1.280 ;
        RECT 2726.750 0.270 2731.150 1.280 ;
        RECT 2732.270 0.270 2736.670 1.280 ;
        RECT 2737.790 0.270 2742.190 1.280 ;
        RECT 2743.310 0.270 2747.710 1.280 ;
        RECT 2748.830 0.270 2753.230 1.280 ;
        RECT 2754.350 0.270 2758.750 1.280 ;
        RECT 2759.870 0.270 2764.270 1.280 ;
        RECT 2765.390 0.270 2769.790 1.280 ;
        RECT 2770.910 0.270 2775.310 1.280 ;
        RECT 2776.430 0.270 2780.830 1.280 ;
        RECT 2781.950 0.270 2786.350 1.280 ;
        RECT 2787.470 0.270 2791.870 1.280 ;
        RECT 2792.990 0.270 2797.390 1.280 ;
        RECT 2798.510 0.270 2870.770 1.280 ;
      LAYER met3 ;
        RECT 1.000 3431.260 2879.000 3468.165 ;
        RECT 1.000 3429.260 2878.600 3431.260 ;
        RECT 1.000 3427.860 2879.000 3429.260 ;
        RECT 1.400 3425.860 2879.000 3427.860 ;
        RECT 1.000 3354.420 2879.000 3425.860 ;
        RECT 1.000 3352.420 2878.600 3354.420 ;
        RECT 1.000 3345.580 2879.000 3352.420 ;
        RECT 1.400 3343.580 2879.000 3345.580 ;
        RECT 1.000 3277.580 2879.000 3343.580 ;
        RECT 1.000 3275.580 2878.600 3277.580 ;
        RECT 1.000 3263.300 2879.000 3275.580 ;
        RECT 1.400 3261.300 2879.000 3263.300 ;
        RECT 1.000 3200.740 2879.000 3261.300 ;
        RECT 1.000 3198.740 2878.600 3200.740 ;
        RECT 1.000 3181.020 2879.000 3198.740 ;
        RECT 1.400 3179.020 2879.000 3181.020 ;
        RECT 1.000 3123.900 2879.000 3179.020 ;
        RECT 1.000 3121.900 2878.600 3123.900 ;
        RECT 1.000 3098.740 2879.000 3121.900 ;
        RECT 1.400 3096.740 2879.000 3098.740 ;
        RECT 1.000 3047.060 2879.000 3096.740 ;
        RECT 1.000 3045.060 2878.600 3047.060 ;
        RECT 1.000 3016.460 2879.000 3045.060 ;
        RECT 1.400 3014.460 2879.000 3016.460 ;
        RECT 1.000 2970.220 2879.000 3014.460 ;
        RECT 1.000 2968.220 2878.600 2970.220 ;
        RECT 1.000 2934.180 2879.000 2968.220 ;
        RECT 1.400 2932.180 2879.000 2934.180 ;
        RECT 1.000 2893.380 2879.000 2932.180 ;
        RECT 1.000 2891.380 2878.600 2893.380 ;
        RECT 1.000 2851.900 2879.000 2891.380 ;
        RECT 1.400 2849.900 2879.000 2851.900 ;
        RECT 1.000 2816.540 2879.000 2849.900 ;
        RECT 1.000 2814.540 2878.600 2816.540 ;
        RECT 1.000 2769.620 2879.000 2814.540 ;
        RECT 1.400 2767.620 2879.000 2769.620 ;
        RECT 1.000 2739.700 2879.000 2767.620 ;
        RECT 1.000 2737.700 2878.600 2739.700 ;
        RECT 1.000 2687.340 2879.000 2737.700 ;
        RECT 1.400 2685.340 2879.000 2687.340 ;
        RECT 1.000 2662.860 2879.000 2685.340 ;
        RECT 1.000 2660.860 2878.600 2662.860 ;
        RECT 1.000 2605.060 2879.000 2660.860 ;
        RECT 1.400 2603.060 2879.000 2605.060 ;
        RECT 1.000 2586.020 2879.000 2603.060 ;
        RECT 1.000 2584.020 2878.600 2586.020 ;
        RECT 1.000 2522.780 2879.000 2584.020 ;
        RECT 1.400 2520.780 2879.000 2522.780 ;
        RECT 1.000 2509.180 2879.000 2520.780 ;
        RECT 1.000 2507.180 2878.600 2509.180 ;
        RECT 1.000 2440.500 2879.000 2507.180 ;
        RECT 1.400 2438.500 2879.000 2440.500 ;
        RECT 1.000 2432.340 2879.000 2438.500 ;
        RECT 1.000 2430.340 2878.600 2432.340 ;
        RECT 1.000 2358.220 2879.000 2430.340 ;
        RECT 1.400 2356.220 2879.000 2358.220 ;
        RECT 1.000 2355.500 2879.000 2356.220 ;
        RECT 1.000 2353.500 2878.600 2355.500 ;
        RECT 1.000 2278.660 2879.000 2353.500 ;
        RECT 1.000 2276.660 2878.600 2278.660 ;
        RECT 1.000 2275.940 2879.000 2276.660 ;
        RECT 1.400 2273.940 2879.000 2275.940 ;
        RECT 1.000 2201.820 2879.000 2273.940 ;
        RECT 1.000 2199.820 2878.600 2201.820 ;
        RECT 1.000 2193.660 2879.000 2199.820 ;
        RECT 1.400 2191.660 2879.000 2193.660 ;
        RECT 1.000 2124.980 2879.000 2191.660 ;
        RECT 1.000 2122.980 2878.600 2124.980 ;
        RECT 1.000 2111.380 2879.000 2122.980 ;
        RECT 1.400 2109.380 2879.000 2111.380 ;
        RECT 1.000 2048.140 2879.000 2109.380 ;
        RECT 1.000 2046.140 2878.600 2048.140 ;
        RECT 1.000 2029.100 2879.000 2046.140 ;
        RECT 1.400 2027.100 2879.000 2029.100 ;
        RECT 1.000 1971.300 2879.000 2027.100 ;
        RECT 1.000 1969.300 2878.600 1971.300 ;
        RECT 1.000 1946.820 2879.000 1969.300 ;
        RECT 1.400 1944.820 2879.000 1946.820 ;
        RECT 1.000 1894.460 2879.000 1944.820 ;
        RECT 1.000 1892.460 2878.600 1894.460 ;
        RECT 1.000 1864.540 2879.000 1892.460 ;
        RECT 1.400 1862.540 2879.000 1864.540 ;
        RECT 1.000 1817.620 2879.000 1862.540 ;
        RECT 1.000 1815.620 2878.600 1817.620 ;
        RECT 1.000 1782.260 2879.000 1815.620 ;
        RECT 1.400 1780.260 2879.000 1782.260 ;
        RECT 1.000 1740.780 2879.000 1780.260 ;
        RECT 1.000 1738.780 2878.600 1740.780 ;
        RECT 1.000 1699.980 2879.000 1738.780 ;
        RECT 1.400 1697.980 2879.000 1699.980 ;
        RECT 1.000 1663.940 2879.000 1697.980 ;
        RECT 1.000 1661.940 2878.600 1663.940 ;
        RECT 1.000 1617.700 2879.000 1661.940 ;
        RECT 1.400 1615.700 2879.000 1617.700 ;
        RECT 1.000 1587.100 2879.000 1615.700 ;
        RECT 1.000 1585.100 2878.600 1587.100 ;
        RECT 1.000 1535.420 2879.000 1585.100 ;
        RECT 1.400 1533.420 2879.000 1535.420 ;
        RECT 1.000 1510.260 2879.000 1533.420 ;
        RECT 1.000 1508.260 2878.600 1510.260 ;
        RECT 1.000 1453.140 2879.000 1508.260 ;
        RECT 1.400 1451.140 2879.000 1453.140 ;
        RECT 1.000 1433.420 2879.000 1451.140 ;
        RECT 1.000 1431.420 2878.600 1433.420 ;
        RECT 1.000 1370.860 2879.000 1431.420 ;
        RECT 1.400 1368.860 2879.000 1370.860 ;
        RECT 1.000 1356.580 2879.000 1368.860 ;
        RECT 1.000 1354.580 2878.600 1356.580 ;
        RECT 1.000 1288.580 2879.000 1354.580 ;
        RECT 1.400 1286.580 2879.000 1288.580 ;
        RECT 1.000 1279.740 2879.000 1286.580 ;
        RECT 1.000 1277.740 2878.600 1279.740 ;
        RECT 1.000 1206.300 2879.000 1277.740 ;
        RECT 1.400 1204.300 2879.000 1206.300 ;
        RECT 1.000 1202.900 2879.000 1204.300 ;
        RECT 1.000 1200.900 2878.600 1202.900 ;
        RECT 1.000 1126.060 2879.000 1200.900 ;
        RECT 1.000 1124.060 2878.600 1126.060 ;
        RECT 1.000 1124.020 2879.000 1124.060 ;
        RECT 1.400 1122.020 2879.000 1124.020 ;
        RECT 1.000 1049.220 2879.000 1122.020 ;
        RECT 1.000 1047.220 2878.600 1049.220 ;
        RECT 1.000 1041.740 2879.000 1047.220 ;
        RECT 1.400 1039.740 2879.000 1041.740 ;
        RECT 1.000 972.380 2879.000 1039.740 ;
        RECT 1.000 970.380 2878.600 972.380 ;
        RECT 1.000 959.460 2879.000 970.380 ;
        RECT 1.400 957.460 2879.000 959.460 ;
        RECT 1.000 895.540 2879.000 957.460 ;
        RECT 1.000 893.540 2878.600 895.540 ;
        RECT 1.000 877.180 2879.000 893.540 ;
        RECT 1.400 875.180 2879.000 877.180 ;
        RECT 1.000 818.700 2879.000 875.180 ;
        RECT 1.000 816.700 2878.600 818.700 ;
        RECT 1.000 794.900 2879.000 816.700 ;
        RECT 1.400 792.900 2879.000 794.900 ;
        RECT 1.000 741.860 2879.000 792.900 ;
        RECT 1.000 739.860 2878.600 741.860 ;
        RECT 1.000 712.620 2879.000 739.860 ;
        RECT 1.400 710.620 2879.000 712.620 ;
        RECT 1.000 665.020 2879.000 710.620 ;
        RECT 1.000 663.020 2878.600 665.020 ;
        RECT 1.000 630.340 2879.000 663.020 ;
        RECT 1.400 628.340 2879.000 630.340 ;
        RECT 1.000 588.180 2879.000 628.340 ;
        RECT 1.000 586.180 2878.600 588.180 ;
        RECT 1.000 548.060 2879.000 586.180 ;
        RECT 1.400 546.060 2879.000 548.060 ;
        RECT 1.000 511.340 2879.000 546.060 ;
        RECT 1.000 509.340 2878.600 511.340 ;
        RECT 1.000 465.780 2879.000 509.340 ;
        RECT 1.400 463.780 2879.000 465.780 ;
        RECT 1.000 434.500 2879.000 463.780 ;
        RECT 1.000 432.500 2878.600 434.500 ;
        RECT 1.000 383.500 2879.000 432.500 ;
        RECT 1.400 381.500 2879.000 383.500 ;
        RECT 1.000 357.660 2879.000 381.500 ;
        RECT 1.000 355.660 2878.600 357.660 ;
        RECT 1.000 301.220 2879.000 355.660 ;
        RECT 1.400 299.220 2879.000 301.220 ;
        RECT 1.000 280.820 2879.000 299.220 ;
        RECT 1.000 278.820 2878.600 280.820 ;
        RECT 1.000 218.940 2879.000 278.820 ;
        RECT 1.400 216.940 2879.000 218.940 ;
        RECT 1.000 203.980 2879.000 216.940 ;
        RECT 1.000 201.980 2878.600 203.980 ;
        RECT 1.000 136.660 2879.000 201.980 ;
        RECT 1.400 134.660 2879.000 136.660 ;
        RECT 1.000 127.140 2879.000 134.660 ;
        RECT 1.000 125.140 2878.600 127.140 ;
        RECT 1.000 54.380 2879.000 125.140 ;
        RECT 1.400 52.380 2879.000 54.380 ;
        RECT 1.000 50.300 2879.000 52.380 ;
        RECT 1.000 48.300 2878.600 50.300 ;
        RECT 1.000 10.715 2879.000 48.300 ;
      LAYER met4 ;
        RECT 7.655 12.415 8.570 3467.145 ;
        RECT 12.470 3378.880 98.570 3467.145 ;
        RECT 12.470 2936.960 45.430 3378.880 ;
        RECT 49.330 3376.140 98.570 3378.880 ;
        RECT 102.470 3376.140 188.570 3467.145 ;
        RECT 192.470 3376.140 278.570 3467.145 ;
        RECT 282.470 3376.140 368.570 3467.145 ;
        RECT 372.470 3376.140 458.570 3467.145 ;
        RECT 462.470 3376.140 548.570 3467.145 ;
        RECT 552.470 3376.140 638.570 3467.145 ;
        RECT 642.470 3376.140 728.570 3467.145 ;
        RECT 732.470 3376.140 818.570 3467.145 ;
        RECT 49.330 2940.400 818.570 3376.140 ;
        RECT 49.330 2936.960 98.570 2940.400 ;
        RECT 12.470 2818.560 98.570 2936.960 ;
        RECT 12.470 2376.640 45.430 2818.560 ;
        RECT 49.330 2816.140 98.570 2818.560 ;
        RECT 102.470 2816.140 188.570 2940.400 ;
        RECT 192.470 2816.140 278.570 2940.400 ;
        RECT 282.470 2816.140 368.570 2940.400 ;
        RECT 372.470 2816.140 458.570 2940.400 ;
        RECT 462.470 2816.140 548.570 2940.400 ;
        RECT 552.470 2816.140 638.570 2940.400 ;
        RECT 642.470 2816.140 728.570 2940.400 ;
        RECT 732.470 2816.140 818.570 2940.400 ;
        RECT 49.330 2380.400 818.570 2816.140 ;
        RECT 49.330 2376.640 98.570 2380.400 ;
        RECT 12.470 2258.240 98.570 2376.640 ;
        RECT 12.470 1816.320 45.430 2258.240 ;
        RECT 49.330 2256.140 98.570 2258.240 ;
        RECT 102.470 2256.140 188.570 2380.400 ;
        RECT 192.470 2256.140 278.570 2380.400 ;
        RECT 282.470 2256.140 368.570 2380.400 ;
        RECT 372.470 2256.140 458.570 2380.400 ;
        RECT 462.470 2256.140 548.570 2380.400 ;
        RECT 552.470 2256.140 638.570 2380.400 ;
        RECT 642.470 2256.140 728.570 2380.400 ;
        RECT 732.470 2256.140 818.570 2380.400 ;
        RECT 49.330 1820.400 818.570 2256.140 ;
        RECT 49.330 1816.320 98.570 1820.400 ;
        RECT 12.470 1697.920 98.570 1816.320 ;
        RECT 12.470 1256.000 45.430 1697.920 ;
        RECT 49.330 1696.140 98.570 1697.920 ;
        RECT 102.470 1696.140 188.570 1820.400 ;
        RECT 192.470 1696.140 278.570 1820.400 ;
        RECT 282.470 1696.140 368.570 1820.400 ;
        RECT 372.470 1696.140 458.570 1820.400 ;
        RECT 462.470 1696.140 548.570 1820.400 ;
        RECT 552.470 1696.140 638.570 1820.400 ;
        RECT 642.470 1696.140 728.570 1820.400 ;
        RECT 732.470 1696.140 818.570 1820.400 ;
        RECT 49.330 1260.400 818.570 1696.140 ;
        RECT 49.330 1256.000 98.570 1260.400 ;
        RECT 12.470 12.415 98.570 1256.000 ;
        RECT 102.470 12.415 188.570 1260.400 ;
        RECT 192.470 12.415 278.570 1260.400 ;
        RECT 282.470 12.415 368.570 1260.400 ;
        RECT 372.470 12.415 458.570 1260.400 ;
        RECT 462.470 12.415 548.570 1260.400 ;
        RECT 552.470 12.415 638.570 1260.400 ;
        RECT 642.470 12.415 728.570 1260.400 ;
        RECT 732.470 12.415 818.570 1260.400 ;
        RECT 822.470 3359.840 908.570 3467.145 ;
        RECT 822.470 2934.240 844.910 3359.840 ;
        RECT 848.810 3357.100 908.570 3359.840 ;
        RECT 912.470 3357.100 998.570 3467.145 ;
        RECT 1002.470 3357.100 1088.570 3467.145 ;
        RECT 1092.470 3357.100 1178.570 3467.145 ;
        RECT 1182.470 3357.100 1268.570 3467.145 ;
        RECT 1272.470 3357.100 1358.570 3467.145 ;
        RECT 1362.470 3362.560 1448.570 3467.145 ;
        RECT 1362.470 3357.100 1437.390 3362.560 ;
        RECT 848.810 2940.400 1437.390 3357.100 ;
        RECT 848.810 2934.240 908.570 2940.400 ;
        RECT 822.470 12.415 908.570 2934.240 ;
        RECT 912.470 12.415 998.570 2940.400 ;
        RECT 1002.470 12.415 1088.570 2940.400 ;
        RECT 1092.470 12.415 1178.570 2940.400 ;
        RECT 1182.470 12.415 1268.570 2940.400 ;
        RECT 1272.470 12.415 1358.570 2940.400 ;
        RECT 1362.470 2936.960 1437.390 2940.400 ;
        RECT 1441.290 2936.960 1448.570 3362.560 ;
        RECT 1362.470 12.415 1448.570 2936.960 ;
        RECT 1452.470 3357.100 1538.570 3467.145 ;
        RECT 1542.470 3357.100 1628.570 3467.145 ;
        RECT 1632.470 3357.100 1718.570 3467.145 ;
        RECT 1722.470 3357.100 1808.570 3467.145 ;
        RECT 1812.470 3357.100 1898.570 3467.145 ;
        RECT 1902.470 3357.100 1988.570 3467.145 ;
        RECT 1452.470 2940.400 1988.570 3357.100 ;
        RECT 1452.470 557.100 1538.570 2940.400 ;
        RECT 1542.470 557.100 1628.570 2940.400 ;
        RECT 1632.470 557.100 1718.570 2940.400 ;
        RECT 1722.470 557.100 1808.570 2940.400 ;
        RECT 1812.470 557.100 1898.570 2940.400 ;
        RECT 1902.470 557.100 1988.570 2940.400 ;
        RECT 1452.470 140.400 1988.570 557.100 ;
        RECT 1452.470 12.415 1538.570 140.400 ;
        RECT 1542.470 12.415 1628.570 140.400 ;
        RECT 1632.470 12.415 1718.570 140.400 ;
        RECT 1722.470 12.415 1808.570 140.400 ;
        RECT 1812.470 12.415 1898.570 140.400 ;
        RECT 1902.470 12.415 1988.570 140.400 ;
        RECT 1992.470 12.415 2078.570 3467.145 ;
        RECT 2082.470 3376.140 2168.570 3467.145 ;
        RECT 2172.470 3376.140 2258.570 3467.145 ;
        RECT 2262.470 3376.140 2348.570 3467.145 ;
        RECT 2352.470 3376.140 2438.570 3467.145 ;
        RECT 2442.470 3376.140 2528.570 3467.145 ;
        RECT 2532.470 3376.140 2618.570 3467.145 ;
        RECT 2622.470 3376.140 2708.570 3467.145 ;
        RECT 2712.470 3376.140 2798.570 3467.145 ;
        RECT 2082.470 2940.400 2798.570 3376.140 ;
        RECT 2082.470 2816.140 2168.570 2940.400 ;
        RECT 2172.470 2816.140 2258.570 2940.400 ;
        RECT 2262.470 2816.140 2348.570 2940.400 ;
        RECT 2352.470 2816.140 2438.570 2940.400 ;
        RECT 2442.470 2816.140 2528.570 2940.400 ;
        RECT 2532.470 2816.140 2618.570 2940.400 ;
        RECT 2622.470 2816.140 2708.570 2940.400 ;
        RECT 2712.470 2816.140 2798.570 2940.400 ;
        RECT 2082.470 2380.400 2798.570 2816.140 ;
        RECT 2082.470 2256.140 2168.570 2380.400 ;
        RECT 2172.470 2256.140 2258.570 2380.400 ;
        RECT 2262.470 2256.140 2348.570 2380.400 ;
        RECT 2352.470 2256.140 2438.570 2380.400 ;
        RECT 2442.470 2256.140 2528.570 2380.400 ;
        RECT 2532.470 2256.140 2618.570 2380.400 ;
        RECT 2622.470 2256.140 2708.570 2380.400 ;
        RECT 2712.470 2256.140 2798.570 2380.400 ;
        RECT 2082.470 1820.400 2798.570 2256.140 ;
        RECT 2082.470 1696.140 2168.570 1820.400 ;
        RECT 2172.470 1696.140 2258.570 1820.400 ;
        RECT 2262.470 1696.140 2348.570 1820.400 ;
        RECT 2352.470 1696.140 2438.570 1820.400 ;
        RECT 2442.470 1696.140 2528.570 1820.400 ;
        RECT 2532.470 1696.140 2618.570 1820.400 ;
        RECT 2622.470 1696.140 2708.570 1820.400 ;
        RECT 2712.470 1696.140 2798.570 1820.400 ;
        RECT 2082.470 1260.400 2798.570 1696.140 ;
        RECT 2082.470 1136.140 2168.570 1260.400 ;
        RECT 2172.470 1136.140 2258.570 1260.400 ;
        RECT 2262.470 1136.140 2348.570 1260.400 ;
        RECT 2352.470 1136.140 2438.570 1260.400 ;
        RECT 2442.470 1136.140 2528.570 1260.400 ;
        RECT 2532.470 1136.140 2618.570 1260.400 ;
        RECT 2622.470 1136.140 2708.570 1260.400 ;
        RECT 2712.470 1136.140 2798.570 1260.400 ;
        RECT 2082.470 700.400 2798.570 1136.140 ;
        RECT 2082.470 576.140 2168.570 700.400 ;
        RECT 2172.470 576.140 2258.570 700.400 ;
        RECT 2262.470 576.140 2348.570 700.400 ;
        RECT 2352.470 576.140 2438.570 700.400 ;
        RECT 2442.470 576.140 2528.570 700.400 ;
        RECT 2532.470 576.140 2618.570 700.400 ;
        RECT 2622.470 576.140 2708.570 700.400 ;
        RECT 2712.470 576.140 2798.570 700.400 ;
        RECT 2082.470 140.400 2798.570 576.140 ;
        RECT 2082.470 12.415 2168.570 140.400 ;
        RECT 2172.470 12.415 2258.570 140.400 ;
        RECT 2262.470 12.415 2348.570 140.400 ;
        RECT 2352.470 12.415 2438.570 140.400 ;
        RECT 2442.470 12.415 2528.570 140.400 ;
        RECT 2532.470 12.415 2618.570 140.400 ;
        RECT 2622.470 12.415 2708.570 140.400 ;
        RECT 2712.470 12.415 2798.570 140.400 ;
        RECT 2802.470 3381.600 2870.530 3467.145 ;
        RECT 2802.470 2934.240 2831.190 3381.600 ;
        RECT 2835.090 2934.240 2870.530 3381.600 ;
        RECT 2802.470 2821.280 2870.530 2934.240 ;
        RECT 2802.470 2379.360 2831.190 2821.280 ;
        RECT 2835.090 2379.360 2870.530 2821.280 ;
        RECT 2802.470 2260.960 2870.530 2379.360 ;
        RECT 2802.470 1819.040 2831.190 2260.960 ;
        RECT 2835.090 1819.040 2870.530 2260.960 ;
        RECT 2802.470 1700.640 2870.530 1819.040 ;
        RECT 2802.470 1258.720 2831.190 1700.640 ;
        RECT 2835.090 1258.720 2870.530 1700.640 ;
        RECT 2802.470 1140.320 2870.530 1258.720 ;
        RECT 2802.470 698.400 2831.190 1140.320 ;
        RECT 2835.090 698.400 2870.530 1140.320 ;
        RECT 2802.470 580.000 2870.530 698.400 ;
        RECT 2802.470 138.080 2831.190 580.000 ;
        RECT 2835.090 138.080 2870.530 580.000 ;
        RECT 2802.470 12.415 2870.530 138.080 ;
      LAYER met5 ;
        RECT 88.900 3079.030 2870.740 3113.500 ;
        RECT 88.900 2989.030 2870.740 3072.730 ;
        RECT 88.900 2899.030 2870.740 2982.730 ;
        RECT 88.900 2881.250 2870.740 2892.730 ;
        RECT 823.670 2874.950 2077.370 2881.250 ;
        RECT 2803.670 2874.950 2870.740 2881.250 ;
        RECT 88.900 2809.030 2870.740 2874.950 ;
        RECT 88.900 2719.030 2870.740 2802.730 ;
        RECT 88.900 2629.030 2870.740 2712.730 ;
        RECT 88.900 2539.030 2870.740 2622.730 ;
        RECT 88.900 2449.030 2870.740 2532.730 ;
        RECT 88.900 2359.030 2870.740 2442.730 ;
        RECT 88.900 2269.030 2870.740 2352.730 ;
        RECT 88.900 2179.030 2870.740 2262.730 ;
        RECT 88.900 2089.030 2870.740 2172.730 ;
        RECT 88.900 1999.030 2870.740 2082.730 ;
        RECT 88.900 1909.030 2870.740 1992.730 ;
        RECT 88.900 1819.030 2870.740 1902.730 ;
        RECT 88.900 1729.030 2870.740 1812.730 ;
        RECT 88.900 1639.030 2870.740 1722.730 ;
        RECT 88.900 1549.030 2870.740 1632.730 ;
        RECT 88.900 1459.030 2870.740 1542.730 ;
        RECT 88.900 1369.030 2870.740 1452.730 ;
        RECT 88.900 1279.030 2870.740 1362.730 ;
        RECT 88.900 1201.650 2870.740 1272.730 ;
        RECT 88.900 1195.350 1987.370 1201.650 ;
        RECT 88.900 1189.030 2870.740 1195.350 ;
        RECT 88.900 1099.030 2870.740 1182.730 ;
        RECT 88.900 1009.030 2870.740 1092.730 ;
        RECT 88.900 919.030 2870.740 1002.730 ;
        RECT 88.900 829.030 2870.740 912.730 ;
        RECT 88.900 739.030 2870.740 822.730 ;
        RECT 88.900 649.030 2870.740 732.730 ;
        RECT 88.900 640.650 2870.740 642.730 ;
        RECT 88.900 634.350 1987.370 640.650 ;
        RECT 88.900 559.030 2870.740 634.350 ;
        RECT 88.900 469.030 2870.740 552.730 ;
        RECT 88.900 379.030 2870.740 462.730 ;
        RECT 88.900 289.030 2870.740 372.730 ;
        RECT 88.900 199.030 2870.740 282.730 ;
        RECT 88.900 140.300 2870.740 192.730 ;
  END
END Marmot
END LIBRARY

