magic
tech sky130B
magscale 1 2
timestamp 1662180296
<< metal1 >>
rect 186498 702992 186504 703044
rect 186556 703032 186562 703044
rect 188430 703032 188436 703044
rect 186556 703004 188436 703032
rect 186556 702992 186562 703004
rect 188430 702992 188436 703004
rect 188488 702992 188494 703044
rect 235166 702992 235172 703044
rect 235224 703032 235230 703044
rect 236178 703032 236184 703044
rect 235224 703004 236184 703032
rect 235224 702992 235230 703004
rect 236178 702992 236184 703004
rect 236236 702992 236242 703044
rect 522758 702992 522764 703044
rect 522816 703032 522822 703044
rect 527082 703032 527088 703044
rect 522816 703004 527088 703032
rect 522816 702992 522822 703004
rect 527082 702992 527088 703004
rect 527140 702992 527146 703044
rect 570506 702992 570512 703044
rect 570564 703032 570570 703044
rect 575842 703032 575848 703044
rect 570564 703004 575848 703032
rect 570564 702992 570570 703004
rect 575842 702992 575848 703004
rect 575900 702992 575906 703044
rect 490926 702720 490932 702772
rect 490984 702760 490990 702772
rect 494790 702760 494796 702772
rect 490984 702732 494796 702760
rect 490984 702720 490990 702732
rect 494790 702720 494796 702732
rect 494848 702720 494854 702772
rect 538674 702720 538680 702772
rect 538732 702760 538738 702772
rect 543458 702760 543464 702772
rect 538732 702732 543464 702760
rect 538732 702720 538738 702732
rect 543458 702720 543464 702732
rect 543516 702720 543522 702772
rect 24302 702448 24308 702500
rect 24360 702488 24366 702500
rect 29270 702488 29276 702500
rect 24360 702460 29276 702488
rect 24360 702448 24366 702460
rect 29270 702448 29276 702460
rect 29328 702448 29334 702500
rect 218974 702448 218980 702500
rect 219032 702488 219038 702500
rect 220262 702488 220268 702500
rect 219032 702460 220268 702488
rect 219032 702448 219038 702460
rect 220262 702448 220268 702460
rect 220320 702448 220326 702500
rect 459094 702448 459100 702500
rect 459152 702488 459158 702500
rect 462314 702488 462320 702500
rect 459152 702460 462320 702488
rect 459152 702448 459158 702460
rect 462314 702448 462320 702460
rect 462372 702448 462378 702500
rect 506842 702448 506848 702500
rect 506900 702488 506906 702500
rect 510982 702488 510988 702500
rect 506900 702460 510988 702488
rect 506900 702448 506906 702460
rect 510982 702448 510988 702460
rect 511040 702448 511046 702500
rect 554590 702448 554596 702500
rect 554648 702488 554654 702500
rect 559650 702488 559656 702500
rect 554648 702460 559656 702488
rect 554648 702448 554654 702460
rect 559650 702448 559656 702460
rect 559708 702448 559714 702500
rect 8110 700952 8116 701004
rect 8168 700992 8174 701004
rect 13078 700992 13084 701004
rect 8168 700964 13084 700992
rect 8168 700952 8174 700964
rect 13078 700952 13084 700964
rect 13136 700952 13142 701004
rect 40494 700952 40500 701004
rect 40552 700992 40558 701004
rect 44910 700992 44916 701004
rect 40552 700964 44916 700992
rect 40552 700952 40558 700964
rect 44910 700952 44916 700964
rect 44968 700952 44974 701004
rect 56778 700952 56784 701004
rect 56836 700992 56842 701004
rect 60734 700992 60740 701004
rect 56836 700964 60740 700992
rect 56836 700952 56842 700964
rect 60734 700952 60740 700964
rect 60792 700952 60798 701004
rect 72970 700952 72976 701004
rect 73028 700992 73034 701004
rect 76742 700992 76748 701004
rect 73028 700964 76748 700992
rect 73028 700952 73034 700964
rect 76742 700952 76748 700964
rect 76800 700952 76806 701004
rect 89162 700952 89168 701004
rect 89220 700992 89226 701004
rect 92566 700992 92572 701004
rect 89220 700964 92572 700992
rect 89220 700952 89226 700964
rect 92566 700952 92572 700964
rect 92624 700952 92630 701004
rect 105446 700952 105452 701004
rect 105504 700992 105510 701004
rect 108574 700992 108580 701004
rect 105504 700964 108580 700992
rect 105504 700952 105510 700964
rect 108574 700952 108580 700964
rect 108632 700952 108638 701004
rect 121638 700952 121644 701004
rect 121696 700992 121702 701004
rect 124398 700992 124404 701004
rect 121696 700964 124404 700992
rect 121696 700952 121702 700964
rect 124398 700952 124404 700964
rect 124456 700952 124462 701004
rect 137830 700952 137836 701004
rect 137888 700992 137894 701004
rect 140406 700992 140412 701004
rect 137888 700964 140412 700992
rect 137888 700952 137894 700964
rect 140406 700952 140412 700964
rect 140464 700952 140470 701004
rect 154114 700952 154120 701004
rect 154172 700992 154178 701004
rect 156230 700992 156236 701004
rect 154172 700964 156236 700992
rect 154172 700952 154178 700964
rect 156230 700952 156236 700964
rect 156288 700952 156294 701004
rect 170306 700952 170312 701004
rect 170364 700992 170370 701004
rect 172422 700992 172428 701004
rect 170364 700964 172428 700992
rect 170364 700952 170370 700964
rect 172422 700952 172428 700964
rect 172480 700952 172486 701004
rect 202782 700952 202788 701004
rect 202840 700992 202846 701004
rect 204254 700992 204260 701004
rect 202840 700964 204260 700992
rect 202840 700952 202846 700964
rect 204254 700952 204260 700964
rect 204312 700952 204318 701004
rect 348050 700952 348056 701004
rect 348108 700992 348114 701004
rect 348786 700992 348792 701004
rect 348108 700964 348792 700992
rect 348108 700952 348114 700964
rect 348786 700952 348792 700964
rect 348844 700952 348850 701004
rect 363874 700952 363880 701004
rect 363932 700992 363938 701004
rect 364978 700992 364984 701004
rect 363932 700964 364984 700992
rect 363932 700952 363938 700964
rect 364978 700952 364984 700964
rect 365036 700952 365042 701004
rect 379330 700952 379336 701004
rect 379388 700992 379394 701004
rect 381170 700992 381176 701004
rect 379388 700964 381176 700992
rect 379388 700952 379394 700964
rect 381170 700952 381176 700964
rect 381228 700952 381234 701004
rect 395706 700952 395712 701004
rect 395764 700992 395770 701004
rect 397454 700992 397460 701004
rect 395764 700964 397460 700992
rect 395764 700952 395770 700964
rect 397454 700952 397460 700964
rect 397512 700952 397518 701004
rect 411714 700952 411720 701004
rect 411772 700992 411778 701004
rect 413646 700992 413652 701004
rect 411772 700964 413652 700992
rect 411772 700952 411778 700964
rect 413646 700952 413652 700964
rect 413704 700952 413710 701004
rect 427538 700952 427544 701004
rect 427596 700992 427602 701004
rect 429838 700992 429844 701004
rect 427596 700964 429844 700992
rect 427596 700952 427602 700964
rect 429838 700952 429844 700964
rect 429896 700952 429902 701004
rect 443546 700952 443552 701004
rect 443604 700992 443610 701004
rect 446122 700992 446128 701004
rect 443604 700964 446128 700992
rect 443604 700952 443610 700964
rect 446122 700952 446128 700964
rect 446180 700952 446186 701004
rect 475378 700952 475384 701004
rect 475436 700992 475442 701004
rect 478506 700992 478512 701004
rect 475436 700964 478512 700992
rect 475436 700952 475442 700964
rect 478506 700952 478512 700964
rect 478564 700952 478570 701004
rect 65518 3816 65524 3868
rect 65576 3856 65582 3868
rect 80238 3856 80244 3868
rect 65576 3828 80244 3856
rect 65576 3816 65582 3828
rect 80238 3816 80244 3828
rect 80296 3816 80302 3868
rect 97626 3816 97632 3868
rect 97684 3856 97690 3868
rect 101214 3856 101220 3868
rect 97684 3828 101220 3856
rect 97684 3816 97690 3828
rect 101214 3816 101220 3828
rect 101272 3816 101278 3868
rect 56042 3748 56048 3800
rect 56100 3788 56106 3800
rect 71406 3788 71412 3800
rect 56100 3760 71412 3788
rect 56100 3748 56106 3760
rect 71406 3748 71412 3760
rect 71464 3748 71470 3800
rect 90082 3748 90088 3800
rect 90140 3788 90146 3800
rect 103422 3788 103428 3800
rect 90140 3760 103428 3788
rect 90140 3748 90146 3760
rect 103422 3748 103428 3760
rect 103480 3748 103486 3800
rect 104342 3748 104348 3800
rect 104400 3788 104406 3800
rect 104400 3760 113174 3788
rect 104400 3748 104406 3760
rect 52546 3680 52552 3732
rect 52604 3720 52610 3732
rect 68094 3720 68100 3732
rect 52604 3692 68100 3720
rect 52604 3680 52610 3692
rect 68094 3680 68100 3692
rect 68152 3680 68158 3732
rect 71866 3680 71872 3732
rect 71924 3720 71930 3732
rect 85758 3720 85764 3732
rect 71924 3692 85764 3720
rect 71924 3680 71930 3692
rect 85758 3680 85764 3692
rect 85816 3680 85822 3732
rect 86862 3680 86868 3732
rect 86920 3720 86926 3732
rect 100110 3720 100116 3732
rect 86920 3692 100116 3720
rect 86920 3680 86926 3692
rect 100110 3680 100116 3692
rect 100168 3680 100174 3732
rect 106642 3680 106648 3732
rect 106700 3720 106706 3732
rect 113146 3720 113174 3760
rect 116670 3720 116676 3732
rect 106700 3692 110184 3720
rect 113146 3692 116676 3720
rect 106700 3680 106706 3692
rect 48958 3612 48964 3664
rect 49016 3652 49022 3664
rect 64782 3652 64788 3664
rect 49016 3624 64788 3652
rect 49016 3612 49022 3624
rect 64782 3612 64788 3624
rect 64840 3612 64846 3664
rect 66714 3612 66720 3664
rect 66772 3652 66778 3664
rect 81434 3652 81440 3664
rect 66772 3624 81440 3652
rect 66772 3612 66778 3624
rect 81434 3612 81440 3624
rect 81492 3612 81498 3664
rect 84470 3612 84476 3664
rect 84528 3652 84534 3664
rect 97902 3652 97908 3664
rect 84528 3624 97908 3652
rect 84528 3612 84534 3624
rect 97902 3612 97908 3624
rect 97960 3612 97966 3664
rect 110046 3652 110052 3664
rect 98012 3624 110052 3652
rect 60826 3544 60832 3596
rect 60884 3584 60890 3596
rect 75914 3584 75920 3596
rect 60884 3556 75920 3584
rect 60884 3544 60890 3556
rect 75914 3544 75920 3556
rect 75972 3544 75978 3596
rect 76282 3544 76288 3596
rect 76340 3584 76346 3596
rect 90174 3584 90180 3596
rect 76340 3556 90180 3584
rect 76340 3544 76346 3556
rect 90174 3544 90180 3556
rect 90232 3544 90238 3596
rect 97626 3584 97632 3596
rect 93826 3556 97632 3584
rect 54938 3476 54944 3528
rect 54996 3516 55002 3528
rect 70302 3516 70308 3528
rect 54996 3488 70308 3516
rect 54996 3476 55002 3488
rect 70302 3476 70308 3488
rect 70360 3476 70366 3528
rect 71498 3476 71504 3528
rect 71556 3516 71562 3528
rect 71866 3516 71872 3528
rect 71556 3488 71872 3516
rect 71556 3476 71562 3488
rect 71866 3476 71872 3488
rect 71924 3476 71930 3528
rect 72970 3476 72976 3528
rect 73028 3516 73034 3528
rect 86954 3516 86960 3528
rect 73028 3488 86960 3516
rect 73028 3476 73034 3488
rect 86954 3476 86960 3488
rect 87012 3476 87018 3528
rect 87782 3476 87788 3528
rect 87840 3516 87846 3528
rect 93826 3516 93854 3556
rect 97626 3544 97632 3556
rect 97684 3544 97690 3596
rect 87840 3488 93854 3516
rect 87840 3476 87846 3488
rect 97442 3476 97448 3528
rect 97500 3516 97506 3528
rect 98012 3516 98040 3624
rect 110046 3612 110052 3624
rect 110104 3612 110110 3664
rect 110156 3652 110184 3692
rect 116670 3680 116676 3692
rect 116728 3680 116734 3732
rect 118878 3652 118884 3664
rect 110156 3624 118884 3652
rect 118878 3612 118884 3624
rect 118936 3612 118942 3664
rect 125962 3612 125968 3664
rect 126020 3652 126026 3664
rect 136542 3652 136548 3664
rect 126020 3624 136548 3652
rect 126020 3612 126026 3624
rect 136542 3612 136548 3624
rect 136600 3612 136606 3664
rect 143626 3612 143632 3664
rect 143684 3652 143690 3664
rect 153194 3652 153200 3664
rect 143684 3624 153200 3652
rect 143684 3612 143690 3624
rect 153194 3612 153200 3624
rect 153252 3612 153258 3664
rect 108482 3544 108488 3596
rect 108540 3584 108546 3596
rect 119982 3584 119988 3596
rect 108540 3556 119988 3584
rect 108540 3544 108546 3556
rect 119982 3544 119988 3556
rect 120040 3544 120046 3596
rect 122282 3544 122288 3596
rect 122340 3584 122346 3596
rect 133230 3584 133236 3596
rect 122340 3556 133236 3584
rect 122340 3544 122346 3556
rect 133230 3544 133236 3556
rect 133288 3544 133294 3596
rect 142522 3544 142528 3596
rect 142580 3584 142586 3596
rect 151998 3584 152004 3596
rect 142580 3556 152004 3584
rect 142580 3544 142586 3556
rect 151998 3544 152004 3556
rect 152056 3544 152062 3596
rect 97500 3488 98040 3516
rect 97500 3476 97506 3488
rect 98638 3476 98644 3528
rect 98696 3516 98702 3528
rect 98696 3488 102456 3516
rect 98696 3476 98702 3488
rect 51350 3408 51356 3460
rect 51408 3448 51414 3460
rect 66990 3448 66996 3460
rect 51408 3420 66996 3448
rect 51408 3408 51414 3420
rect 66990 3408 66996 3420
rect 67048 3408 67054 3460
rect 70118 3408 70124 3460
rect 70176 3448 70182 3460
rect 84654 3448 84660 3460
rect 70176 3420 84660 3448
rect 70176 3408 70182 3420
rect 84654 3408 84660 3420
rect 84712 3408 84718 3460
rect 89530 3408 89536 3460
rect 89588 3448 89594 3460
rect 102318 3448 102324 3460
rect 89588 3420 102324 3448
rect 89588 3408 89594 3420
rect 102318 3408 102324 3420
rect 102376 3408 102382 3460
rect 102428 3448 102456 3488
rect 110506 3476 110512 3528
rect 110564 3516 110570 3528
rect 122374 3516 122380 3528
rect 110564 3488 122380 3516
rect 110564 3476 110570 3488
rect 122374 3476 122380 3488
rect 122432 3476 122438 3528
rect 129366 3476 129372 3528
rect 129424 3516 129430 3528
rect 139854 3516 139860 3528
rect 129424 3488 139860 3516
rect 129424 3476 129430 3488
rect 139854 3476 139860 3488
rect 139912 3476 139918 3528
rect 141602 3476 141608 3528
rect 141660 3516 141666 3528
rect 150894 3516 150900 3528
rect 141660 3488 150900 3516
rect 141660 3476 141666 3488
rect 150894 3476 150900 3488
rect 150952 3476 150958 3528
rect 111150 3448 111156 3460
rect 102428 3420 111156 3448
rect 111150 3408 111156 3420
rect 111208 3408 111214 3460
rect 117590 3408 117596 3460
rect 117648 3448 117654 3460
rect 128814 3448 128820 3460
rect 117648 3420 128820 3448
rect 117648 3408 117654 3420
rect 128814 3408 128820 3420
rect 128872 3408 128878 3460
rect 138750 3448 138756 3460
rect 128924 3420 138756 3448
rect 63218 3340 63224 3392
rect 63276 3380 63282 3392
rect 78030 3380 78036 3392
rect 63276 3352 78036 3380
rect 63276 3340 63282 3352
rect 78030 3340 78036 3352
rect 78088 3340 78094 3392
rect 83274 3340 83280 3392
rect 83332 3380 83338 3392
rect 92934 3380 92940 3392
rect 83332 3352 92940 3380
rect 83332 3340 83338 3352
rect 92934 3340 92940 3352
rect 92992 3340 92998 3392
rect 93946 3340 93952 3392
rect 94004 3380 94010 3392
rect 94004 3352 99512 3380
rect 94004 3340 94010 3352
rect 62022 3272 62028 3324
rect 62080 3312 62086 3324
rect 76926 3312 76932 3324
rect 62080 3284 76932 3312
rect 62080 3272 62086 3284
rect 76926 3272 76932 3284
rect 76984 3272 76990 3324
rect 82078 3272 82084 3324
rect 82136 3312 82142 3324
rect 95694 3312 95700 3324
rect 82136 3284 95700 3312
rect 82136 3272 82142 3284
rect 95694 3272 95700 3284
rect 95752 3272 95758 3324
rect 58802 3204 58808 3256
rect 58860 3244 58866 3256
rect 73614 3244 73620 3256
rect 58860 3216 73620 3244
rect 58860 3204 58866 3216
rect 73614 3204 73620 3216
rect 73672 3204 73678 3256
rect 77386 3204 77392 3256
rect 77444 3244 77450 3256
rect 91278 3244 91284 3256
rect 77444 3216 91284 3244
rect 77444 3204 77450 3216
rect 91278 3204 91284 3216
rect 91336 3204 91342 3256
rect 96246 3204 96252 3256
rect 96304 3244 96310 3256
rect 99484 3244 99512 3352
rect 101030 3340 101036 3392
rect 101088 3380 101094 3392
rect 113358 3380 113364 3392
rect 101088 3352 113364 3380
rect 101088 3340 101094 3352
rect 113358 3340 113364 3352
rect 113416 3340 113422 3392
rect 116394 3340 116400 3392
rect 116452 3380 116458 3392
rect 121546 3380 121552 3392
rect 116452 3352 121552 3380
rect 116452 3340 116458 3352
rect 121546 3340 121552 3352
rect 121604 3340 121610 3392
rect 128170 3340 128176 3392
rect 128228 3380 128234 3392
rect 128924 3380 128952 3420
rect 138750 3408 138756 3420
rect 138808 3408 138814 3460
rect 149790 3448 149796 3460
rect 141068 3420 149796 3448
rect 128228 3352 128952 3380
rect 128228 3340 128234 3352
rect 130562 3340 130568 3392
rect 130620 3380 130626 3392
rect 140682 3380 140688 3392
rect 130620 3352 140688 3380
rect 130620 3340 130626 3352
rect 140682 3340 140688 3352
rect 140740 3340 140746 3392
rect 103330 3272 103336 3324
rect 103388 3312 103394 3324
rect 115566 3312 115572 3324
rect 103388 3284 115572 3312
rect 103388 3272 103394 3284
rect 115566 3272 115572 3284
rect 115624 3272 115630 3324
rect 119890 3272 119896 3324
rect 119948 3312 119954 3324
rect 131022 3312 131028 3324
rect 119948 3284 131028 3312
rect 119948 3272 119954 3284
rect 131022 3272 131028 3284
rect 131080 3272 131086 3324
rect 140038 3272 140044 3324
rect 140096 3312 140102 3324
rect 141068 3312 141096 3420
rect 149790 3408 149796 3420
rect 149848 3408 149854 3460
rect 147582 3380 147588 3392
rect 140096 3284 141096 3312
rect 141160 3352 147588 3380
rect 140096 3272 140102 3284
rect 106734 3244 106740 3256
rect 96304 3216 99420 3244
rect 99484 3216 106740 3244
rect 96304 3204 96310 3216
rect 56962 3136 56968 3188
rect 57020 3176 57026 3188
rect 72510 3176 72516 3188
rect 57020 3148 72516 3176
rect 57020 3136 57026 3148
rect 72510 3136 72516 3148
rect 72568 3136 72574 3188
rect 73798 3136 73804 3188
rect 73856 3176 73862 3188
rect 87966 3176 87972 3188
rect 73856 3148 87972 3176
rect 73856 3136 73862 3148
rect 87966 3136 87972 3148
rect 88024 3136 88030 3188
rect 92842 3136 92848 3188
rect 92900 3176 92906 3188
rect 99392 3176 99420 3216
rect 106734 3204 106740 3216
rect 106792 3204 106798 3256
rect 111610 3204 111616 3256
rect 111668 3244 111674 3256
rect 123294 3244 123300 3256
rect 111668 3216 123300 3244
rect 111668 3204 111674 3216
rect 123294 3204 123300 3216
rect 123352 3204 123358 3256
rect 123754 3204 123760 3256
rect 123812 3244 123818 3256
rect 134334 3244 134340 3256
rect 123812 3216 134340 3244
rect 123812 3204 123818 3216
rect 134334 3204 134340 3216
rect 134392 3204 134398 3256
rect 137646 3204 137652 3256
rect 137704 3244 137710 3256
rect 141160 3244 141188 3352
rect 147582 3340 147588 3352
rect 147640 3340 147646 3392
rect 154022 3340 154028 3392
rect 154080 3380 154086 3392
rect 163038 3380 163044 3392
rect 154080 3352 163044 3380
rect 154080 3340 154086 3352
rect 163038 3340 163044 3352
rect 163096 3340 163102 3392
rect 166074 3340 166080 3392
rect 166132 3380 166138 3392
rect 174078 3380 174084 3392
rect 166132 3352 174084 3380
rect 166132 3340 166138 3352
rect 174078 3340 174084 3352
rect 174136 3340 174142 3392
rect 183738 3340 183744 3392
rect 183796 3380 183802 3392
rect 190638 3380 190644 3392
rect 183796 3352 190644 3380
rect 183796 3340 183802 3352
rect 190638 3340 190644 3352
rect 190696 3340 190702 3392
rect 553302 3340 553308 3392
rect 553360 3380 553366 3392
rect 571518 3380 571524 3392
rect 553360 3352 571524 3380
rect 553360 3340 553366 3352
rect 571518 3340 571524 3352
rect 571576 3340 571582 3392
rect 145926 3272 145932 3324
rect 145984 3312 145990 3324
rect 155310 3312 155316 3324
rect 145984 3284 155316 3312
rect 145984 3272 145990 3284
rect 155310 3272 155316 3284
rect 155368 3272 155374 3324
rect 155770 3272 155776 3324
rect 155828 3312 155834 3324
rect 164234 3312 164240 3324
rect 155828 3284 164240 3312
rect 155828 3272 155834 3284
rect 164234 3272 164240 3284
rect 164292 3272 164298 3324
rect 164878 3272 164884 3324
rect 164936 3312 164942 3324
rect 172974 3312 172980 3324
rect 164936 3284 172980 3312
rect 164936 3272 164942 3284
rect 172974 3272 172980 3284
rect 173032 3272 173038 3324
rect 176746 3272 176752 3324
rect 176804 3312 176810 3324
rect 184014 3312 184020 3324
rect 176804 3284 184020 3312
rect 176804 3272 176810 3284
rect 184014 3272 184020 3284
rect 184072 3272 184078 3324
rect 184934 3272 184940 3324
rect 184992 3312 184998 3324
rect 184992 3284 190454 3312
rect 184992 3272 184998 3284
rect 137704 3216 141188 3244
rect 137704 3204 137710 3216
rect 151814 3204 151820 3256
rect 151872 3244 151878 3256
rect 160830 3244 160836 3256
rect 151872 3216 160836 3244
rect 151872 3204 151878 3216
rect 160830 3204 160836 3216
rect 160888 3204 160894 3256
rect 162486 3204 162492 3256
rect 162544 3244 162550 3256
rect 170766 3244 170772 3256
rect 162544 3216 170772 3244
rect 162544 3204 162550 3216
rect 170766 3204 170772 3216
rect 170824 3204 170830 3256
rect 171870 3244 171876 3256
rect 171106 3216 171876 3244
rect 108942 3176 108948 3188
rect 92900 3148 98684 3176
rect 99392 3148 108948 3176
rect 92900 3136 92906 3148
rect 40954 3068 40960 3120
rect 41012 3108 41018 3120
rect 57054 3108 57060 3120
rect 41012 3080 57060 3108
rect 41012 3068 41018 3080
rect 57054 3068 57060 3080
rect 57112 3068 57118 3120
rect 80882 3068 80888 3120
rect 80940 3108 80946 3120
rect 94590 3108 94596 3120
rect 80940 3080 94596 3108
rect 80940 3068 80946 3080
rect 94590 3068 94596 3080
rect 94648 3068 94654 3120
rect 98656 3108 98684 3148
rect 108942 3136 108948 3148
rect 109000 3136 109006 3188
rect 109402 3136 109408 3188
rect 109460 3176 109466 3188
rect 121086 3176 121092 3188
rect 109460 3148 121092 3176
rect 109460 3136 109466 3148
rect 121086 3136 121092 3148
rect 121144 3136 121150 3188
rect 132126 3176 132132 3188
rect 121196 3148 132132 3176
rect 121196 3120 121224 3148
rect 132126 3136 132132 3148
rect 132184 3136 132190 3188
rect 136450 3136 136456 3188
rect 136508 3176 136514 3188
rect 146202 3176 146208 3188
rect 136508 3148 146208 3176
rect 136508 3136 136514 3148
rect 146202 3136 146208 3148
rect 146260 3136 146266 3188
rect 154206 3176 154212 3188
rect 146312 3148 154212 3176
rect 105630 3108 105636 3120
rect 98656 3080 105636 3108
rect 105630 3068 105636 3080
rect 105688 3068 105694 3120
rect 106090 3068 106096 3120
rect 106148 3108 106154 3120
rect 117774 3108 117780 3120
rect 106148 3080 117780 3108
rect 106148 3068 106154 3080
rect 117774 3068 117780 3080
rect 117832 3068 117838 3120
rect 121178 3068 121184 3120
rect 121236 3068 121242 3120
rect 121546 3068 121552 3120
rect 121604 3108 121610 3120
rect 127710 3108 127716 3120
rect 121604 3080 127716 3108
rect 121604 3068 121610 3080
rect 127710 3068 127716 3080
rect 127768 3068 127774 3120
rect 131758 3068 131764 3120
rect 131816 3108 131822 3120
rect 142062 3108 142068 3120
rect 131816 3080 142068 3108
rect 131816 3068 131822 3080
rect 142062 3068 142068 3080
rect 142120 3068 142126 3120
rect 144730 3068 144736 3120
rect 144788 3108 144794 3120
rect 146312 3108 146340 3148
rect 154206 3136 154212 3148
rect 154264 3136 154270 3188
rect 156322 3136 156328 3188
rect 156380 3176 156386 3188
rect 165246 3176 165252 3188
rect 156380 3148 165252 3176
rect 156380 3136 156386 3148
rect 165246 3136 165252 3148
rect 165304 3136 165310 3188
rect 165706 3136 165712 3188
rect 165764 3176 165770 3188
rect 171106 3176 171134 3216
rect 171870 3204 171876 3216
rect 171928 3204 171934 3256
rect 173158 3204 173164 3256
rect 173216 3244 173222 3256
rect 180886 3244 180892 3256
rect 173216 3216 180892 3244
rect 173216 3204 173222 3216
rect 180886 3204 180892 3216
rect 180944 3204 180950 3256
rect 181438 3204 181444 3256
rect 181496 3244 181502 3256
rect 188430 3244 188436 3256
rect 181496 3216 188436 3244
rect 181496 3204 181502 3216
rect 188430 3204 188436 3216
rect 188488 3204 188494 3256
rect 190426 3244 190454 3284
rect 550082 3272 550088 3324
rect 550140 3312 550146 3324
rect 568022 3312 568028 3324
rect 550140 3284 568028 3312
rect 550140 3272 550146 3284
rect 568022 3272 568028 3284
rect 568080 3272 568086 3324
rect 191834 3244 191840 3256
rect 190426 3216 191840 3244
rect 191834 3204 191840 3216
rect 191892 3204 191898 3256
rect 197354 3244 197360 3256
rect 194244 3216 197360 3244
rect 165764 3148 171134 3176
rect 165764 3136 165770 3148
rect 174262 3136 174268 3188
rect 174320 3176 174326 3188
rect 174320 3148 176424 3176
rect 174320 3136 174326 3148
rect 144788 3080 146340 3108
rect 144788 3068 144794 3080
rect 149514 3068 149520 3120
rect 149572 3108 149578 3120
rect 158714 3108 158720 3120
rect 149572 3080 158720 3108
rect 149572 3068 149578 3080
rect 158714 3068 158720 3080
rect 158772 3068 158778 3120
rect 160186 3068 160192 3120
rect 160244 3108 160250 3120
rect 168558 3108 168564 3120
rect 160244 3080 168564 3108
rect 160244 3068 160250 3080
rect 168558 3068 168564 3080
rect 168616 3068 168622 3120
rect 176286 3108 176292 3120
rect 168668 3080 176292 3108
rect 50154 3000 50160 3052
rect 50212 3040 50218 3052
rect 65886 3040 65892 3052
rect 50212 3012 65892 3040
rect 50212 3000 50218 3012
rect 65886 3000 65892 3012
rect 65944 3000 65950 3052
rect 69106 3000 69112 3052
rect 69164 3040 69170 3052
rect 83550 3040 83556 3052
rect 69164 3012 83556 3040
rect 69164 3000 69170 3012
rect 83550 3000 83556 3012
rect 83608 3000 83614 3052
rect 92382 3040 92388 3052
rect 84166 3012 92388 3040
rect 26602 2932 26608 2984
rect 26660 2972 26666 2984
rect 44082 2972 44088 2984
rect 26660 2944 44088 2972
rect 26660 2932 26666 2944
rect 44082 2932 44088 2944
rect 44140 2932 44146 2984
rect 44266 2932 44272 2984
rect 44324 2972 44330 2984
rect 44324 2944 45554 2972
rect 44324 2932 44330 2944
rect 27706 2864 27712 2916
rect 27764 2904 27770 2916
rect 45186 2904 45192 2916
rect 27764 2876 45192 2904
rect 27764 2864 27770 2876
rect 45186 2864 45192 2876
rect 45244 2864 45250 2916
rect 45526 2904 45554 2944
rect 47854 2932 47860 2984
rect 47912 2972 47918 2984
rect 63402 2972 63408 2984
rect 47912 2944 63408 2972
rect 47912 2932 47918 2944
rect 63402 2932 63408 2944
rect 63460 2932 63466 2984
rect 67910 2932 67916 2984
rect 67968 2972 67974 2984
rect 77110 2972 77116 2984
rect 67968 2944 77116 2972
rect 67968 2932 67974 2944
rect 77110 2932 77116 2944
rect 77168 2932 77174 2984
rect 78582 2932 78588 2984
rect 78640 2972 78646 2984
rect 84166 2972 84194 3012
rect 92382 3000 92388 3012
rect 92440 3000 92446 3052
rect 95142 3040 95148 3052
rect 92584 3012 95148 3040
rect 88978 2972 88984 2984
rect 78640 2944 84194 2972
rect 85592 2944 88984 2972
rect 78640 2932 78646 2944
rect 60642 2904 60648 2916
rect 45526 2876 60648 2904
rect 60642 2864 60648 2876
rect 60700 2864 60706 2916
rect 74994 2904 75000 2916
rect 60844 2876 75000 2904
rect 33594 2796 33600 2848
rect 33652 2836 33658 2848
rect 50706 2836 50712 2848
rect 33652 2808 50712 2836
rect 33652 2796 33658 2808
rect 50706 2796 50712 2808
rect 50764 2796 50770 2848
rect 59630 2796 59636 2848
rect 59688 2836 59694 2848
rect 60844 2836 60872 2876
rect 74994 2864 75000 2876
rect 75052 2864 75058 2916
rect 75362 2864 75368 2916
rect 75420 2904 75426 2916
rect 85482 2904 85488 2916
rect 75420 2876 85488 2904
rect 75420 2864 75426 2876
rect 85482 2864 85488 2876
rect 85540 2864 85546 2916
rect 59688 2808 60872 2836
rect 59688 2796 59694 2808
rect 64322 2796 64328 2848
rect 64380 2836 64386 2848
rect 68830 2836 68836 2848
rect 64380 2808 68836 2836
rect 64380 2796 64386 2808
rect 68830 2796 68836 2808
rect 68888 2796 68894 2848
rect 79686 2796 79692 2848
rect 79744 2836 79750 2848
rect 85592 2836 85620 2944
rect 88978 2932 88984 2944
rect 89036 2932 89042 2984
rect 85666 2864 85672 2916
rect 85724 2904 85730 2916
rect 92584 2904 92612 3012
rect 95142 3000 95148 3012
rect 95200 3000 95206 3052
rect 104526 3040 104532 3052
rect 97736 3012 104532 3040
rect 97736 2972 97764 3012
rect 104526 3000 104532 3012
rect 104584 3000 104590 3052
rect 112806 3000 112812 3052
rect 112864 3040 112870 3052
rect 124398 3040 124404 3052
rect 112864 3012 124404 3040
rect 112864 3000 112870 3012
rect 124398 3000 124404 3012
rect 124456 3000 124462 3052
rect 125042 3000 125048 3052
rect 125100 3040 125106 3052
rect 135162 3040 135168 3052
rect 125100 3012 135168 3040
rect 125100 3000 125106 3012
rect 135162 3000 135168 3012
rect 135220 3000 135226 3052
rect 135898 3000 135904 3052
rect 135956 3040 135962 3052
rect 145374 3040 145380 3052
rect 135956 3012 145380 3040
rect 135956 3000 135962 3012
rect 145374 3000 145380 3012
rect 145432 3000 145438 3052
rect 147122 3000 147128 3052
rect 147180 3040 147186 3052
rect 156414 3040 156420 3052
rect 147180 3012 156420 3040
rect 147180 3000 147186 3012
rect 156414 3000 156420 3012
rect 156472 3000 156478 3052
rect 159266 3000 159272 3052
rect 159324 3040 159330 3052
rect 167454 3040 167460 3052
rect 159324 3012 167460 3040
rect 159324 3000 159330 3012
rect 167454 3000 167460 3012
rect 167512 3000 167518 3052
rect 168374 3000 168380 3052
rect 168432 3040 168438 3052
rect 168668 3040 168696 3080
rect 176286 3068 176292 3080
rect 176344 3068 176350 3120
rect 176396 3108 176424 3148
rect 179046 3136 179052 3188
rect 179104 3176 179110 3188
rect 186314 3176 186320 3188
rect 179104 3148 186320 3176
rect 179104 3136 179110 3148
rect 186314 3136 186320 3148
rect 186372 3136 186378 3188
rect 190822 3136 190828 3188
rect 190880 3176 190886 3188
rect 194244 3176 194272 3216
rect 197354 3204 197360 3216
rect 197412 3204 197418 3256
rect 214466 3204 214472 3256
rect 214524 3244 214530 3256
rect 219342 3244 219348 3256
rect 214524 3216 219348 3244
rect 214524 3204 214530 3216
rect 219342 3204 219348 3216
rect 219400 3204 219406 3256
rect 530026 3204 530032 3256
rect 530084 3244 530090 3256
rect 546678 3244 546684 3256
rect 530084 3216 546684 3244
rect 530084 3204 530090 3216
rect 546678 3204 546684 3216
rect 546736 3204 546742 3256
rect 556706 3204 556712 3256
rect 556764 3244 556770 3256
rect 575106 3244 575112 3256
rect 556764 3216 575112 3244
rect 556764 3204 556770 3216
rect 575106 3204 575112 3216
rect 575164 3204 575170 3256
rect 190880 3148 194272 3176
rect 190880 3136 190886 3148
rect 196802 3136 196808 3188
rect 196860 3176 196866 3188
rect 202874 3176 202880 3188
rect 196860 3148 202880 3176
rect 196860 3136 196866 3148
rect 202874 3136 202880 3148
rect 202932 3136 202938 3188
rect 209866 3136 209872 3188
rect 209924 3176 209930 3188
rect 214926 3176 214932 3188
rect 209924 3148 214932 3176
rect 209924 3136 209930 3148
rect 214926 3136 214932 3148
rect 214984 3136 214990 3188
rect 220446 3136 220452 3188
rect 220504 3176 220510 3188
rect 224862 3176 224868 3188
rect 220504 3148 224868 3176
rect 220504 3136 220510 3148
rect 224862 3136 224868 3148
rect 224920 3136 224926 3188
rect 561122 3136 561128 3188
rect 561180 3176 561186 3188
rect 579798 3176 579804 3188
rect 561180 3148 579804 3176
rect 561180 3136 561186 3148
rect 579798 3136 579804 3148
rect 579856 3136 579862 3188
rect 181806 3108 181812 3120
rect 176396 3080 181812 3108
rect 181806 3068 181812 3080
rect 181864 3068 181870 3120
rect 186130 3068 186136 3120
rect 186188 3108 186194 3120
rect 192846 3108 192852 3120
rect 186188 3080 192852 3108
rect 186188 3068 186194 3080
rect 192846 3068 192852 3080
rect 192904 3068 192910 3120
rect 193306 3068 193312 3120
rect 193364 3108 193370 3120
rect 199470 3108 199476 3120
rect 193364 3080 199476 3108
rect 193364 3068 193370 3080
rect 199470 3068 199476 3080
rect 199528 3068 199534 3120
rect 200298 3068 200304 3120
rect 200356 3108 200362 3120
rect 206094 3108 206100 3120
rect 200356 3080 206100 3108
rect 200356 3068 200362 3080
rect 206094 3068 206100 3080
rect 206152 3068 206158 3120
rect 206186 3068 206192 3120
rect 206244 3108 206250 3120
rect 211614 3108 211620 3120
rect 206244 3080 211620 3108
rect 206244 3068 206250 3080
rect 211614 3068 211620 3080
rect 211672 3068 211678 3120
rect 216858 3068 216864 3120
rect 216916 3108 216922 3120
rect 221550 3108 221556 3120
rect 216916 3080 221556 3108
rect 216916 3068 216922 3080
rect 221550 3068 221556 3080
rect 221608 3068 221614 3120
rect 231026 3068 231032 3120
rect 231084 3108 231090 3120
rect 234798 3108 234804 3120
rect 231084 3080 234804 3108
rect 231084 3068 231090 3080
rect 234798 3068 234804 3080
rect 234856 3068 234862 3120
rect 239306 3068 239312 3120
rect 239364 3108 239370 3120
rect 242526 3108 242532 3120
rect 239364 3080 242532 3108
rect 239364 3068 239370 3080
rect 242526 3068 242532 3080
rect 242584 3068 242590 3120
rect 532602 3068 532608 3120
rect 532660 3108 532666 3120
rect 540790 3108 540796 3120
rect 532660 3080 540796 3108
rect 532660 3068 532666 3080
rect 540790 3068 540796 3080
rect 540848 3068 540854 3120
rect 563146 3068 563152 3120
rect 563204 3108 563210 3120
rect 582190 3108 582196 3120
rect 563204 3080 582196 3108
rect 563204 3068 563210 3080
rect 582190 3068 582196 3080
rect 582248 3068 582254 3120
rect 175274 3040 175280 3052
rect 168432 3012 168696 3040
rect 171106 3012 175280 3040
rect 168432 3000 168438 3012
rect 85724 2876 92612 2904
rect 93826 2944 97764 2972
rect 85724 2864 85730 2876
rect 79744 2808 85620 2836
rect 79744 2796 79750 2808
rect 91922 2796 91928 2848
rect 91980 2836 91986 2848
rect 93826 2836 93854 2944
rect 102226 2932 102232 2984
rect 102284 2972 102290 2984
rect 102284 2944 113174 2972
rect 102284 2932 102290 2944
rect 95050 2864 95056 2916
rect 95108 2904 95114 2916
rect 107838 2904 107844 2916
rect 95108 2876 107844 2904
rect 95108 2864 95114 2876
rect 107838 2864 107844 2876
rect 107896 2864 107902 2916
rect 113146 2904 113174 2944
rect 114002 2932 114008 2984
rect 114060 2972 114066 2984
rect 125594 2972 125600 2984
rect 114060 2944 125600 2972
rect 114060 2932 114066 2944
rect 125594 2932 125600 2944
rect 125652 2932 125658 2984
rect 134150 2932 134156 2984
rect 134208 2972 134214 2984
rect 144546 2972 144552 2984
rect 134208 2944 144552 2972
rect 134208 2932 134214 2944
rect 144546 2932 144552 2944
rect 144604 2932 144610 2984
rect 148962 2972 148968 2984
rect 145576 2944 148968 2972
rect 114554 2904 114560 2916
rect 113146 2876 114560 2904
rect 114554 2864 114560 2876
rect 114612 2864 114618 2916
rect 115198 2864 115204 2916
rect 115256 2904 115262 2916
rect 126606 2904 126612 2916
rect 115256 2876 126612 2904
rect 115256 2864 115262 2876
rect 126606 2864 126612 2876
rect 126664 2864 126670 2916
rect 126974 2864 126980 2916
rect 127032 2904 127038 2916
rect 137922 2904 137928 2916
rect 127032 2876 137928 2904
rect 127032 2864 127038 2876
rect 137922 2864 137928 2876
rect 137980 2864 137986 2916
rect 138842 2864 138848 2916
rect 138900 2904 138906 2916
rect 145576 2904 145604 2944
rect 148962 2932 148968 2944
rect 149020 2932 149026 2984
rect 153010 2932 153016 2984
rect 153068 2972 153074 2984
rect 162210 2972 162216 2984
rect 153068 2944 162216 2972
rect 153068 2932 153074 2944
rect 162210 2932 162216 2944
rect 162268 2932 162274 2984
rect 163682 2932 163688 2984
rect 163740 2972 163746 2984
rect 165706 2972 165712 2984
rect 163740 2944 165712 2972
rect 163740 2932 163746 2944
rect 165706 2932 165712 2944
rect 165764 2932 165770 2984
rect 167178 2932 167184 2984
rect 167236 2972 167242 2984
rect 171106 2972 171134 3012
rect 175274 3000 175280 3012
rect 175332 3000 175338 3052
rect 175826 3000 175832 3052
rect 175884 3040 175890 3052
rect 182910 3040 182916 3052
rect 175884 3012 182916 3040
rect 175884 3000 175890 3012
rect 182910 3000 182916 3012
rect 182968 3000 182974 3052
rect 188522 3000 188528 3052
rect 188580 3040 188586 3052
rect 195054 3040 195060 3052
rect 188580 3012 195060 3040
rect 188580 3000 188586 3012
rect 195054 3000 195060 3012
rect 195112 3000 195118 3052
rect 195606 3000 195612 3052
rect 195664 3040 195670 3052
rect 201678 3040 201684 3052
rect 195664 3012 201684 3040
rect 195664 3000 195670 3012
rect 201678 3000 201684 3012
rect 201736 3000 201742 3052
rect 206922 3040 206928 3052
rect 201788 3012 206928 3040
rect 167236 2944 171134 2972
rect 167236 2932 167242 2944
rect 171962 2932 171968 2984
rect 172020 2972 172026 2984
rect 179874 2972 179880 2984
rect 172020 2944 179880 2972
rect 172020 2932 172026 2944
rect 179874 2932 179880 2944
rect 179932 2932 179938 2984
rect 182542 2932 182548 2984
rect 182600 2972 182606 2984
rect 189534 2972 189540 2984
rect 182600 2944 189540 2972
rect 182600 2932 182606 2944
rect 189534 2932 189540 2944
rect 189592 2932 189598 2984
rect 189718 2932 189724 2984
rect 189776 2972 189782 2984
rect 196434 2972 196440 2984
rect 189776 2944 196440 2972
rect 189776 2932 189782 2944
rect 196434 2932 196440 2944
rect 196492 2932 196498 2984
rect 201494 2932 201500 2984
rect 201552 2972 201558 2984
rect 201788 2972 201816 3012
rect 206922 3000 206928 3012
rect 206980 3000 206986 3052
rect 210970 3000 210976 3052
rect 211028 3040 211034 3052
rect 216030 3040 216036 3052
rect 211028 3012 216036 3040
rect 211028 3000 211034 3012
rect 216030 3000 216036 3012
rect 216088 3000 216094 3052
rect 218054 3000 218060 3052
rect 218112 3040 218118 3052
rect 222654 3040 222660 3052
rect 218112 3012 222660 3040
rect 218112 3000 218118 3012
rect 222654 3000 222660 3012
rect 222712 3000 222718 3052
rect 225506 3000 225512 3052
rect 225564 3040 225570 3052
rect 229278 3040 229284 3052
rect 225564 3012 229284 3040
rect 225564 3000 225570 3012
rect 229278 3000 229284 3012
rect 229336 3000 229342 3052
rect 229830 3000 229836 3052
rect 229888 3040 229894 3052
rect 233694 3040 233700 3052
rect 229888 3012 233700 3040
rect 229888 3000 229894 3012
rect 233694 3000 233700 3012
rect 233752 3000 233758 3052
rect 234614 3000 234620 3052
rect 234672 3040 234678 3052
rect 238110 3040 238116 3052
rect 234672 3012 238116 3040
rect 234672 3000 234678 3012
rect 238110 3000 238116 3012
rect 238168 3000 238174 3052
rect 240502 3000 240508 3052
rect 240560 3040 240566 3052
rect 243630 3040 243636 3052
rect 240560 3012 243636 3040
rect 240560 3000 240566 3012
rect 243630 3000 243636 3012
rect 243688 3000 243694 3052
rect 248782 3000 248788 3052
rect 248840 3040 248846 3052
rect 251358 3040 251364 3052
rect 248840 3012 251364 3040
rect 248840 3000 248846 3012
rect 251358 3000 251364 3012
rect 251416 3000 251422 3052
rect 331306 3000 331312 3052
rect 331364 3040 331370 3052
rect 333882 3040 333888 3052
rect 331364 3012 333888 3040
rect 331364 3000 331370 3012
rect 333882 3000 333888 3012
rect 333940 3000 333946 3052
rect 334802 3000 334808 3052
rect 334860 3040 334866 3052
rect 337470 3040 337476 3052
rect 334860 3012 337476 3040
rect 334860 3000 334866 3012
rect 337470 3000 337476 3012
rect 337528 3000 337534 3052
rect 513466 3000 513472 3052
rect 513524 3040 513530 3052
rect 529014 3040 529020 3052
rect 513524 3012 529020 3040
rect 513524 3000 513530 3012
rect 529014 3000 529020 3012
rect 529072 3000 529078 3052
rect 535546 3000 535552 3052
rect 535604 3040 535610 3052
rect 542814 3040 542820 3052
rect 535604 3012 542820 3040
rect 535604 3000 535610 3012
rect 542814 3000 542820 3012
rect 542872 3000 542878 3052
rect 543458 3000 543464 3052
rect 543516 3040 543522 3052
rect 560478 3040 560484 3052
rect 543516 3012 560484 3040
rect 543516 3000 543522 3012
rect 560478 3000 560484 3012
rect 560536 3000 560542 3052
rect 564342 3000 564348 3052
rect 564400 3040 564406 3052
rect 583386 3040 583392 3052
rect 564400 3012 583392 3040
rect 564400 3000 564406 3012
rect 583386 3000 583392 3012
rect 583444 3000 583450 3052
rect 201552 2944 201816 2972
rect 201552 2932 201558 2944
rect 203886 2932 203892 2984
rect 203944 2972 203950 2984
rect 209406 2972 209412 2984
rect 203944 2944 209412 2972
rect 203944 2932 203950 2944
rect 209406 2932 209412 2944
rect 209464 2932 209470 2984
rect 212166 2932 212172 2984
rect 212224 2972 212230 2984
rect 217134 2972 217140 2984
rect 212224 2944 217140 2972
rect 212224 2932 212230 2944
rect 217134 2932 217140 2944
rect 217192 2932 217198 2984
rect 222746 2932 222752 2984
rect 222804 2972 222810 2984
rect 227346 2972 227352 2984
rect 222804 2944 227352 2972
rect 222804 2932 222810 2944
rect 227346 2932 227352 2944
rect 227404 2932 227410 2984
rect 227530 2932 227536 2984
rect 227588 2972 227594 2984
rect 231762 2972 231768 2984
rect 227588 2944 231768 2972
rect 227588 2932 227594 2944
rect 231762 2932 231768 2944
rect 231820 2932 231826 2984
rect 232222 2932 232228 2984
rect 232280 2972 232286 2984
rect 236178 2972 236184 2984
rect 232280 2944 236184 2972
rect 232280 2932 232286 2944
rect 236178 2932 236184 2944
rect 236236 2932 236242 2984
rect 237006 2932 237012 2984
rect 237064 2972 237070 2984
rect 240594 2972 240600 2984
rect 237064 2944 240600 2972
rect 237064 2932 237070 2944
rect 240594 2932 240600 2944
rect 240652 2932 240658 2984
rect 242894 2932 242900 2984
rect 242952 2972 242958 2984
rect 246114 2972 246120 2984
rect 242952 2944 246120 2972
rect 242952 2932 242958 2944
rect 246114 2932 246120 2944
rect 246172 2932 246178 2984
rect 246390 2932 246396 2984
rect 246448 2972 246454 2984
rect 249426 2972 249432 2984
rect 246448 2944 249432 2972
rect 246448 2932 246454 2944
rect 249426 2932 249432 2944
rect 249484 2932 249490 2984
rect 253474 2932 253480 2984
rect 253532 2972 253538 2984
rect 256050 2972 256056 2984
rect 253532 2944 256056 2972
rect 253532 2932 253538 2944
rect 256050 2932 256056 2944
rect 256108 2932 256114 2984
rect 310238 2932 310244 2984
rect 310296 2972 310302 2984
rect 311434 2972 311440 2984
rect 310296 2944 311440 2972
rect 310296 2932 310302 2944
rect 311434 2932 311440 2944
rect 311492 2932 311498 2984
rect 325694 2932 325700 2984
rect 325752 2972 325758 2984
rect 327994 2972 328000 2984
rect 325752 2944 328000 2972
rect 325752 2932 325758 2944
rect 327994 2932 328000 2944
rect 328052 2932 328058 2984
rect 329006 2932 329012 2984
rect 329064 2972 329070 2984
rect 331582 2972 331588 2984
rect 329064 2944 331588 2972
rect 329064 2932 329070 2944
rect 331582 2932 331588 2944
rect 331640 2932 331646 2984
rect 332318 2932 332324 2984
rect 332376 2972 332382 2984
rect 335078 2972 335084 2984
rect 332376 2944 335084 2972
rect 332376 2932 332382 2944
rect 335078 2932 335084 2944
rect 335136 2932 335142 2984
rect 341150 2932 341156 2984
rect 341208 2972 341214 2984
rect 344554 2972 344560 2984
rect 341208 2944 344560 2972
rect 341208 2932 341214 2944
rect 344554 2932 344560 2944
rect 344612 2932 344618 2984
rect 514846 2932 514852 2984
rect 514904 2972 514910 2984
rect 521838 2972 521844 2984
rect 514904 2944 521844 2972
rect 514904 2932 514910 2944
rect 521838 2932 521844 2944
rect 521896 2932 521902 2984
rect 536558 2932 536564 2984
rect 536616 2972 536622 2984
rect 553762 2972 553768 2984
rect 536616 2944 553768 2972
rect 536616 2932 536622 2944
rect 553762 2932 553768 2944
rect 553820 2932 553826 2984
rect 138900 2876 145604 2904
rect 138900 2864 138906 2876
rect 148318 2864 148324 2916
rect 148376 2904 148382 2916
rect 157518 2904 157524 2916
rect 148376 2876 157524 2904
rect 148376 2864 148382 2876
rect 157518 2864 157524 2876
rect 157576 2864 157582 2916
rect 157794 2864 157800 2916
rect 157852 2904 157858 2916
rect 166626 2904 166632 2916
rect 157852 2876 166632 2904
rect 157852 2864 157858 2876
rect 166626 2864 166632 2876
rect 166684 2864 166690 2916
rect 169570 2864 169576 2916
rect 169628 2904 169634 2916
rect 177666 2904 177672 2916
rect 169628 2876 177672 2904
rect 169628 2864 169634 2876
rect 177666 2864 177672 2876
rect 177724 2864 177730 2916
rect 177850 2864 177856 2916
rect 177908 2904 177914 2916
rect 185394 2904 185400 2916
rect 177908 2876 185400 2904
rect 177908 2864 177914 2876
rect 185394 2864 185400 2876
rect 185452 2864 185458 2916
rect 187602 2904 187608 2916
rect 185504 2876 187608 2904
rect 91980 2808 93854 2836
rect 91980 2796 91986 2808
rect 99834 2796 99840 2848
rect 99892 2836 99898 2848
rect 112254 2836 112260 2848
rect 99892 2808 112260 2836
rect 99892 2796 99898 2808
rect 112254 2796 112260 2808
rect 112312 2796 112318 2848
rect 118786 2796 118792 2848
rect 118844 2836 118850 2848
rect 129642 2836 129648 2848
rect 118844 2808 129648 2836
rect 118844 2796 118850 2808
rect 129642 2796 129648 2808
rect 129700 2796 129706 2848
rect 132954 2796 132960 2848
rect 133012 2836 133018 2848
rect 143442 2836 143448 2848
rect 133012 2808 143448 2836
rect 133012 2796 133018 2808
rect 143442 2796 143448 2808
rect 143500 2796 143506 2848
rect 150618 2796 150624 2848
rect 150676 2836 150682 2848
rect 160002 2836 160008 2848
rect 150676 2808 160008 2836
rect 150676 2796 150682 2808
rect 160002 2796 160008 2808
rect 160060 2796 160066 2848
rect 161290 2796 161296 2848
rect 161348 2836 161354 2848
rect 169938 2836 169944 2848
rect 161348 2808 169944 2836
rect 161348 2796 161354 2808
rect 169938 2796 169944 2808
rect 169996 2796 170002 2848
rect 170766 2796 170772 2848
rect 170824 2836 170830 2848
rect 178770 2836 178776 2848
rect 170824 2808 178776 2836
rect 170824 2796 170830 2808
rect 178770 2796 178776 2808
rect 178828 2796 178834 2848
rect 180242 2796 180248 2848
rect 180300 2836 180306 2848
rect 185504 2836 185532 2876
rect 187602 2864 187608 2876
rect 187660 2864 187666 2916
rect 192386 2864 192392 2916
rect 192444 2904 192450 2916
rect 198366 2904 198372 2916
rect 192444 2876 198372 2904
rect 192444 2864 192450 2876
rect 198366 2864 198372 2876
rect 198424 2864 198430 2916
rect 199102 2864 199108 2916
rect 199160 2904 199166 2916
rect 204990 2904 204996 2916
rect 199160 2876 204996 2904
rect 199160 2864 199166 2876
rect 204990 2864 204996 2876
rect 205048 2864 205054 2916
rect 205082 2864 205088 2916
rect 205140 2904 205146 2916
rect 210510 2904 210516 2916
rect 205140 2876 210516 2904
rect 205140 2864 205146 2876
rect 210510 2864 210516 2876
rect 210568 2864 210574 2916
rect 213362 2864 213368 2916
rect 213420 2904 213426 2916
rect 218238 2904 218244 2916
rect 213420 2876 218244 2904
rect 213420 2864 213426 2876
rect 218238 2864 218244 2876
rect 218296 2864 218302 2916
rect 219250 2864 219256 2916
rect 219308 2904 219314 2916
rect 223482 2904 223488 2916
rect 219308 2876 223488 2904
rect 219308 2864 219314 2876
rect 223482 2864 223488 2876
rect 223540 2864 223546 2916
rect 223942 2864 223948 2916
rect 224000 2904 224006 2916
rect 228450 2904 228456 2916
rect 224000 2876 228456 2904
rect 224000 2864 224006 2876
rect 228450 2864 228456 2876
rect 228508 2864 228514 2916
rect 228726 2864 228732 2916
rect 228784 2904 228790 2916
rect 232866 2904 232872 2916
rect 228784 2876 232872 2904
rect 228784 2864 228790 2876
rect 232866 2864 232872 2876
rect 232924 2864 232930 2916
rect 235810 2864 235816 2916
rect 235868 2904 235874 2916
rect 239490 2904 239496 2916
rect 235868 2876 239496 2904
rect 235868 2864 235874 2876
rect 239490 2864 239496 2876
rect 239548 2864 239554 2916
rect 242066 2864 242072 2916
rect 242124 2904 242130 2916
rect 245010 2904 245016 2916
rect 242124 2876 245016 2904
rect 242124 2864 242130 2876
rect 245010 2864 245016 2876
rect 245068 2864 245074 2916
rect 245194 2864 245200 2916
rect 245252 2904 245258 2916
rect 248322 2904 248328 2916
rect 245252 2876 248328 2904
rect 245252 2864 245258 2876
rect 248322 2864 248328 2876
rect 248380 2864 248386 2916
rect 249978 2864 249984 2916
rect 250036 2904 250042 2916
rect 252738 2904 252744 2916
rect 250036 2876 252744 2904
rect 250036 2864 250042 2876
rect 252738 2864 252744 2876
rect 252796 2864 252802 2916
rect 254670 2864 254676 2916
rect 254728 2904 254734 2916
rect 257154 2904 257160 2916
rect 254728 2876 257160 2904
rect 254728 2864 254734 2876
rect 257154 2864 257160 2876
rect 257212 2864 257218 2916
rect 261754 2864 261760 2916
rect 261812 2904 261818 2916
rect 263778 2904 263784 2916
rect 261812 2876 263784 2904
rect 261812 2864 261818 2876
rect 263778 2864 263784 2876
rect 263836 2864 263842 2916
rect 312446 2864 312452 2916
rect 312504 2904 312510 2916
rect 313826 2904 313832 2916
rect 312504 2876 313832 2904
rect 312504 2864 312510 2876
rect 313826 2864 313832 2876
rect 313884 2864 313890 2916
rect 314562 2864 314568 2916
rect 314620 2904 314626 2916
rect 316218 2904 316224 2916
rect 314620 2876 316224 2904
rect 314620 2864 314626 2876
rect 316218 2864 316224 2876
rect 316276 2864 316282 2916
rect 316862 2864 316868 2916
rect 316920 2904 316926 2916
rect 318518 2904 318524 2916
rect 316920 2876 318524 2904
rect 316920 2864 316926 2876
rect 318518 2864 318524 2876
rect 318576 2864 318582 2916
rect 319070 2864 319076 2916
rect 319128 2904 319134 2916
rect 320910 2904 320916 2916
rect 319128 2876 320916 2904
rect 319128 2864 319134 2876
rect 320910 2864 320916 2876
rect 320968 2864 320974 2916
rect 321278 2864 321284 2916
rect 321336 2904 321342 2916
rect 323302 2904 323308 2916
rect 321336 2876 323308 2904
rect 321336 2864 321342 2876
rect 323302 2864 323308 2876
rect 323360 2864 323366 2916
rect 323486 2864 323492 2916
rect 323544 2904 323550 2916
rect 325602 2904 325608 2916
rect 323544 2876 325608 2904
rect 323544 2864 323550 2876
rect 325602 2864 325608 2876
rect 325660 2864 325666 2916
rect 327902 2864 327908 2916
rect 327960 2904 327966 2916
rect 330386 2904 330392 2916
rect 327960 2876 330392 2904
rect 327960 2864 327966 2876
rect 330386 2864 330392 2876
rect 330444 2864 330450 2916
rect 333422 2864 333428 2916
rect 333480 2904 333486 2916
rect 336274 2904 336280 2916
rect 333480 2876 336280 2904
rect 333480 2864 333486 2876
rect 336274 2864 336280 2876
rect 336332 2864 336338 2916
rect 340046 2864 340052 2916
rect 340104 2904 340110 2916
rect 342990 2904 342996 2916
rect 340104 2876 342996 2904
rect 340104 2864 340110 2876
rect 342990 2864 342996 2876
rect 343048 2864 343054 2916
rect 514754 2864 514760 2916
rect 514812 2904 514818 2916
rect 523034 2904 523040 2916
rect 514812 2876 523040 2904
rect 514812 2864 514818 2876
rect 523034 2864 523040 2876
rect 523092 2864 523098 2916
rect 525794 2864 525800 2916
rect 525852 2904 525858 2916
rect 531314 2904 531320 2916
rect 525852 2876 531320 2904
rect 525852 2864 525858 2876
rect 531314 2864 531320 2876
rect 531372 2864 531378 2916
rect 532234 2864 532240 2916
rect 532292 2904 532298 2916
rect 539594 2904 539600 2916
rect 532292 2876 539600 2904
rect 532292 2864 532298 2876
rect 539594 2864 539600 2876
rect 539652 2864 539658 2916
rect 541986 2904 541992 2916
rect 541452 2876 541992 2904
rect 180300 2808 185532 2836
rect 180300 2796 180306 2808
rect 187326 2796 187332 2848
rect 187384 2836 187390 2848
rect 194226 2836 194232 2848
rect 187384 2808 194232 2836
rect 187384 2796 187390 2808
rect 194226 2796 194232 2808
rect 194284 2796 194290 2848
rect 194410 2796 194416 2848
rect 194468 2836 194474 2848
rect 200850 2836 200856 2848
rect 194468 2808 200856 2836
rect 194468 2796 194474 2808
rect 200850 2796 200856 2808
rect 200908 2796 200914 2848
rect 202690 2796 202696 2848
rect 202748 2836 202754 2848
rect 208394 2836 208400 2848
rect 202748 2808 208400 2836
rect 202748 2796 202754 2808
rect 208394 2796 208400 2808
rect 208452 2796 208458 2848
rect 208578 2796 208584 2848
rect 208636 2836 208642 2848
rect 213822 2836 213828 2848
rect 208636 2808 213828 2836
rect 208636 2796 208642 2808
rect 213822 2796 213828 2808
rect 213880 2796 213886 2848
rect 215662 2796 215668 2848
rect 215720 2836 215726 2848
rect 220722 2836 220728 2848
rect 215720 2808 220728 2836
rect 215720 2796 215726 2808
rect 220722 2796 220728 2808
rect 220780 2796 220786 2848
rect 221550 2796 221556 2848
rect 221608 2836 221614 2848
rect 226242 2836 226248 2848
rect 221608 2808 226248 2836
rect 221608 2796 221614 2808
rect 226242 2796 226248 2808
rect 226300 2796 226306 2848
rect 226334 2796 226340 2848
rect 226392 2836 226398 2848
rect 230658 2836 230664 2848
rect 226392 2808 230664 2836
rect 226392 2796 226398 2808
rect 230658 2796 230664 2808
rect 230716 2796 230722 2848
rect 233418 2796 233424 2848
rect 233476 2836 233482 2848
rect 237282 2836 237288 2848
rect 233476 2808 237288 2836
rect 233476 2796 233482 2808
rect 237282 2796 237288 2808
rect 237340 2796 237346 2848
rect 238110 2796 238116 2848
rect 238168 2836 238174 2848
rect 241698 2836 241704 2848
rect 238168 2808 241704 2836
rect 238168 2796 238174 2808
rect 241698 2796 241704 2808
rect 241756 2796 241762 2848
rect 244090 2796 244096 2848
rect 244148 2836 244154 2848
rect 247218 2836 247224 2848
rect 244148 2808 247224 2836
rect 244148 2796 244154 2808
rect 247218 2796 247224 2808
rect 247276 2796 247282 2848
rect 247586 2796 247592 2848
rect 247644 2836 247650 2848
rect 250530 2836 250536 2848
rect 247644 2808 250536 2836
rect 247644 2796 247650 2808
rect 250530 2796 250536 2808
rect 250588 2796 250594 2848
rect 252370 2796 252376 2848
rect 252428 2836 252434 2848
rect 254946 2836 254952 2848
rect 252428 2808 254952 2836
rect 252428 2796 252434 2808
rect 254946 2796 254952 2808
rect 255004 2796 255010 2848
rect 255866 2796 255872 2848
rect 255924 2836 255930 2848
rect 258258 2836 258264 2848
rect 255924 2808 258264 2836
rect 255924 2796 255930 2808
rect 258258 2796 258264 2808
rect 258316 2796 258322 2848
rect 260650 2796 260656 2848
rect 260708 2836 260714 2848
rect 262674 2836 262680 2848
rect 260708 2808 262680 2836
rect 260708 2796 260714 2808
rect 262674 2796 262680 2808
rect 262732 2796 262738 2848
rect 304718 2796 304724 2848
rect 304776 2836 304782 2848
rect 305546 2836 305552 2848
rect 304776 2808 305552 2836
rect 304776 2796 304782 2808
rect 305546 2796 305552 2808
rect 305604 2796 305610 2848
rect 306926 2796 306932 2848
rect 306984 2836 306990 2848
rect 307938 2836 307944 2848
rect 306984 2808 307944 2836
rect 306984 2796 306990 2808
rect 307938 2796 307944 2808
rect 307996 2796 308002 2848
rect 309134 2796 309140 2848
rect 309192 2836 309198 2848
rect 310238 2836 310244 2848
rect 309192 2808 310244 2836
rect 309192 2796 309198 2808
rect 310238 2796 310244 2808
rect 310296 2796 310302 2848
rect 311342 2796 311348 2848
rect 311400 2836 311406 2848
rect 312630 2836 312636 2848
rect 311400 2808 312636 2836
rect 311400 2796 311406 2808
rect 312630 2796 312636 2808
rect 312688 2796 312694 2848
rect 313550 2796 313556 2848
rect 313608 2836 313614 2848
rect 315022 2836 315028 2848
rect 313608 2808 315028 2836
rect 313608 2796 313614 2808
rect 315022 2796 315028 2808
rect 315080 2796 315086 2848
rect 315758 2796 315764 2848
rect 315816 2836 315822 2848
rect 317322 2836 317328 2848
rect 315816 2808 317328 2836
rect 315816 2796 315822 2808
rect 317322 2796 317328 2808
rect 317380 2796 317386 2848
rect 317966 2796 317972 2848
rect 318024 2836 318030 2848
rect 319714 2836 319720 2848
rect 318024 2808 319720 2836
rect 318024 2796 318030 2808
rect 319714 2796 319720 2808
rect 319772 2796 319778 2848
rect 320082 2796 320088 2848
rect 320140 2836 320146 2848
rect 322106 2836 322112 2848
rect 320140 2808 322112 2836
rect 320140 2796 320146 2808
rect 322106 2796 322112 2808
rect 322164 2796 322170 2848
rect 322382 2796 322388 2848
rect 322440 2836 322446 2848
rect 324406 2836 324412 2848
rect 322440 2808 324412 2836
rect 322440 2796 322446 2808
rect 324406 2796 324412 2808
rect 324464 2796 324470 2848
rect 324590 2796 324596 2848
rect 324648 2836 324654 2848
rect 326798 2836 326804 2848
rect 324648 2808 326804 2836
rect 324648 2796 324654 2808
rect 326798 2796 326804 2808
rect 326856 2796 326862 2848
rect 326982 2796 326988 2848
rect 327040 2836 327046 2848
rect 329190 2836 329196 2848
rect 327040 2808 329196 2836
rect 327040 2796 327046 2808
rect 329190 2796 329196 2808
rect 329248 2796 329254 2848
rect 330110 2796 330116 2848
rect 330168 2836 330174 2848
rect 332686 2836 332692 2848
rect 330168 2808 332692 2836
rect 330168 2796 330174 2808
rect 332686 2796 332692 2808
rect 332744 2796 332750 2848
rect 335630 2796 335636 2848
rect 335688 2836 335694 2848
rect 338666 2836 338672 2848
rect 335688 2808 338672 2836
rect 335688 2796 335694 2808
rect 338666 2796 338672 2808
rect 338724 2796 338730 2848
rect 338942 2796 338948 2848
rect 339000 2836 339006 2848
rect 342070 2836 342076 2848
rect 339000 2808 342076 2836
rect 339000 2796 339006 2808
rect 342070 2796 342076 2808
rect 342128 2796 342134 2848
rect 346670 2796 346676 2848
rect 346728 2836 346734 2848
rect 350442 2836 350448 2848
rect 346728 2808 350448 2836
rect 346728 2796 346734 2808
rect 350442 2796 350448 2808
rect 350500 2796 350506 2848
rect 353202 2796 353208 2848
rect 353260 2836 353266 2848
rect 357526 2836 357532 2848
rect 353260 2808 357532 2836
rect 353260 2796 353266 2808
rect 357526 2796 357532 2808
rect 357584 2796 357590 2848
rect 372338 2796 372344 2848
rect 372396 2836 372402 2848
rect 377674 2836 377680 2848
rect 372396 2808 377680 2836
rect 372396 2796 372402 2808
rect 377674 2796 377680 2808
rect 377732 2796 377738 2848
rect 520182 2796 520188 2848
rect 520240 2836 520246 2848
rect 520240 2808 525472 2836
rect 520240 2796 520246 2808
rect 525444 2780 525472 2808
rect 536834 2796 536840 2848
rect 536892 2836 536898 2848
rect 541452 2836 541480 2876
rect 541986 2864 541992 2876
rect 542044 2864 542050 2916
rect 561950 2864 561956 2916
rect 562008 2904 562014 2916
rect 580994 2904 581000 2916
rect 562008 2876 581000 2904
rect 562008 2864 562014 2876
rect 580994 2864 581000 2876
rect 581052 2864 581058 2916
rect 536892 2808 541480 2836
rect 536892 2796 536898 2808
rect 541526 2796 541532 2848
rect 541584 2836 541590 2848
rect 550266 2836 550272 2848
rect 541584 2808 550272 2836
rect 541584 2796 541590 2808
rect 550266 2796 550272 2808
rect 550324 2796 550330 2848
rect 559742 2796 559748 2848
rect 559800 2836 559806 2848
rect 578602 2836 578608 2848
rect 559800 2808 578608 2836
rect 559800 2796 559806 2808
rect 578602 2796 578608 2808
rect 578660 2796 578666 2848
rect 525426 2728 525432 2780
rect 525484 2728 525490 2780
rect 77110 1300 77116 1352
rect 77168 1340 77174 1352
rect 82722 1340 82728 1352
rect 77168 1312 82728 1340
rect 77168 1300 77174 1312
rect 82722 1300 82728 1312
rect 82780 1300 82786 1352
rect 88978 1300 88984 1352
rect 89036 1340 89042 1352
rect 93762 1340 93768 1352
rect 89036 1312 93768 1340
rect 89036 1300 89042 1312
rect 93762 1300 93768 1312
rect 93820 1300 93826 1352
rect 95142 1300 95148 1352
rect 95200 1340 95206 1352
rect 99282 1340 99288 1352
rect 95200 1312 99288 1340
rect 95200 1300 95206 1312
rect 99282 1300 99288 1312
rect 99340 1300 99346 1352
rect 198274 1300 198280 1352
rect 198332 1340 198338 1352
rect 204162 1340 204168 1352
rect 198332 1312 204168 1340
rect 198332 1300 198338 1312
rect 204162 1300 204168 1312
rect 204220 1300 204226 1352
rect 207382 1300 207388 1352
rect 207440 1340 207446 1352
rect 212994 1340 213000 1352
rect 207440 1312 213000 1340
rect 207440 1300 207446 1312
rect 212994 1300 213000 1312
rect 213052 1300 213058 1352
rect 257062 1300 257068 1352
rect 257120 1340 257126 1352
rect 259362 1340 259368 1352
rect 257120 1312 259368 1340
rect 257120 1300 257126 1312
rect 259362 1300 259368 1312
rect 259420 1300 259426 1352
rect 259454 1300 259460 1352
rect 259512 1340 259518 1352
rect 261570 1340 261576 1352
rect 259512 1312 261576 1340
rect 259512 1300 259518 1312
rect 261570 1300 261576 1312
rect 261628 1300 261634 1352
rect 262950 1300 262956 1352
rect 263008 1340 263014 1352
rect 264882 1340 264888 1352
rect 263008 1312 264888 1340
rect 263008 1300 263014 1312
rect 264882 1300 264888 1312
rect 264940 1300 264946 1352
rect 265342 1300 265348 1352
rect 265400 1340 265406 1352
rect 267090 1340 267096 1352
rect 265400 1312 267096 1340
rect 265400 1300 265406 1312
rect 267090 1300 267096 1312
rect 267148 1300 267154 1352
rect 267734 1300 267740 1352
rect 267792 1340 267798 1352
rect 269298 1340 269304 1352
rect 267792 1312 269304 1340
rect 267792 1300 267798 1312
rect 269298 1300 269304 1312
rect 269356 1300 269362 1352
rect 271230 1300 271236 1352
rect 271288 1340 271294 1352
rect 272610 1340 272616 1352
rect 271288 1312 272616 1340
rect 271288 1300 271294 1312
rect 272610 1300 272616 1312
rect 272668 1300 272674 1352
rect 273622 1300 273628 1352
rect 273680 1340 273686 1352
rect 274818 1340 274824 1352
rect 273680 1312 274824 1340
rect 273680 1300 273686 1312
rect 274818 1300 274824 1312
rect 274876 1300 274882 1352
rect 277118 1300 277124 1352
rect 277176 1340 277182 1352
rect 278130 1340 278136 1352
rect 277176 1312 278136 1340
rect 277176 1300 277182 1312
rect 278130 1300 278136 1312
rect 278188 1300 278194 1352
rect 279510 1300 279516 1352
rect 279568 1340 279574 1352
rect 280338 1340 280344 1352
rect 279568 1312 280344 1340
rect 279568 1300 279574 1312
rect 280338 1300 280344 1312
rect 280396 1300 280402 1352
rect 336642 1300 336648 1352
rect 336700 1340 336706 1352
rect 339862 1340 339868 1352
rect 336700 1312 339868 1340
rect 336700 1300 336706 1312
rect 339862 1300 339868 1312
rect 339920 1300 339926 1352
rect 342162 1300 342168 1352
rect 342220 1340 342226 1352
rect 345750 1340 345756 1352
rect 342220 1312 345756 1340
rect 342220 1300 342226 1312
rect 345750 1300 345756 1312
rect 345808 1300 345814 1352
rect 348878 1300 348884 1352
rect 348936 1340 348942 1352
rect 352834 1340 352840 1352
rect 348936 1312 352840 1340
rect 348936 1300 348942 1312
rect 352834 1300 352840 1312
rect 352892 1300 352898 1352
rect 356606 1300 356612 1352
rect 356664 1340 356670 1352
rect 361114 1340 361120 1352
rect 356664 1312 361120 1340
rect 356664 1300 356670 1312
rect 361114 1300 361120 1312
rect 361172 1300 361178 1352
rect 364242 1300 364248 1352
rect 364300 1340 364306 1352
rect 369394 1340 369400 1352
rect 364300 1312 369400 1340
rect 364300 1300 364306 1312
rect 369394 1300 369400 1312
rect 369452 1300 369458 1352
rect 374270 1300 374276 1352
rect 374328 1340 374334 1352
rect 379606 1340 379612 1352
rect 374328 1312 379612 1340
rect 374328 1300 374334 1312
rect 379606 1300 379612 1312
rect 379664 1300 379670 1352
rect 385310 1300 385316 1352
rect 385368 1340 385374 1352
rect 391842 1340 391848 1352
rect 385368 1312 391848 1340
rect 385368 1300 385374 1312
rect 391842 1300 391848 1312
rect 391900 1300 391906 1352
rect 396350 1300 396356 1352
rect 396408 1340 396414 1352
rect 403618 1340 403624 1352
rect 396408 1312 403624 1340
rect 396408 1300 396414 1312
rect 403618 1300 403624 1312
rect 403676 1300 403682 1352
rect 406286 1300 406292 1352
rect 406344 1340 406350 1352
rect 414290 1340 414296 1352
rect 406344 1312 414296 1340
rect 406344 1300 406350 1312
rect 414290 1300 414296 1312
rect 414348 1300 414354 1352
rect 415118 1300 415124 1352
rect 415176 1340 415182 1352
rect 423398 1340 423404 1352
rect 415176 1312 423404 1340
rect 415176 1300 415182 1312
rect 423398 1300 423404 1312
rect 423456 1300 423462 1352
rect 428366 1300 428372 1352
rect 428424 1340 428430 1352
rect 437566 1340 437572 1352
rect 428424 1312 437572 1340
rect 428424 1300 428430 1312
rect 437566 1300 437572 1312
rect 437624 1300 437630 1352
rect 439406 1300 439412 1352
rect 439464 1340 439470 1352
rect 443730 1340 443736 1352
rect 439464 1312 443736 1340
rect 439464 1300 439470 1312
rect 443730 1300 443736 1312
rect 443788 1300 443794 1352
rect 445846 1340 445852 1352
rect 443840 1312 445852 1340
rect 85482 1232 85488 1284
rect 85540 1272 85546 1284
rect 89346 1272 89352 1284
rect 85540 1244 89352 1272
rect 85540 1232 85546 1244
rect 89346 1232 89352 1244
rect 89404 1232 89410 1284
rect 92934 1232 92940 1284
rect 92992 1272 92998 1284
rect 97074 1272 97080 1284
rect 92992 1244 97080 1272
rect 92992 1232 92998 1244
rect 97074 1232 97080 1244
rect 97132 1232 97138 1284
rect 258258 1232 258264 1284
rect 258316 1272 258322 1284
rect 260466 1272 260472 1284
rect 258316 1244 260472 1272
rect 258316 1232 258322 1244
rect 260466 1232 260472 1244
rect 260524 1232 260530 1284
rect 264146 1232 264152 1284
rect 264204 1272 264210 1284
rect 265986 1272 265992 1284
rect 264204 1244 265992 1272
rect 264204 1232 264210 1244
rect 265986 1232 265992 1244
rect 266044 1232 266050 1284
rect 266538 1232 266544 1284
rect 266596 1272 266602 1284
rect 268194 1272 268200 1284
rect 266596 1244 268200 1272
rect 266596 1232 266602 1244
rect 268194 1232 268200 1244
rect 268252 1232 268258 1284
rect 270034 1232 270040 1284
rect 270092 1272 270098 1284
rect 271506 1272 271512 1284
rect 270092 1244 271512 1272
rect 270092 1232 270098 1244
rect 271506 1232 271512 1244
rect 271564 1232 271570 1284
rect 272426 1232 272432 1284
rect 272484 1272 272490 1284
rect 273714 1272 273720 1284
rect 272484 1244 273720 1272
rect 272484 1232 272490 1244
rect 273714 1232 273720 1244
rect 273772 1232 273778 1284
rect 343358 1232 343364 1284
rect 343416 1272 343422 1284
rect 346946 1272 346952 1284
rect 343416 1244 346952 1272
rect 343416 1232 343422 1244
rect 346946 1232 346952 1244
rect 347004 1232 347010 1284
rect 349982 1232 349988 1284
rect 350040 1272 350046 1284
rect 354030 1272 354036 1284
rect 350040 1244 354036 1272
rect 350040 1232 350046 1244
rect 354030 1232 354036 1244
rect 354088 1232 354094 1284
rect 357710 1232 357716 1284
rect 357768 1272 357774 1284
rect 362310 1272 362316 1284
rect 357768 1244 362316 1272
rect 357768 1232 357774 1244
rect 362310 1232 362316 1244
rect 362368 1232 362374 1284
rect 365438 1232 365444 1284
rect 365496 1272 365502 1284
rect 370222 1272 370228 1284
rect 365496 1244 370228 1272
rect 365496 1232 365502 1244
rect 370222 1232 370228 1244
rect 370280 1232 370286 1284
rect 370958 1232 370964 1284
rect 371016 1272 371022 1284
rect 376110 1272 376116 1284
rect 371016 1244 376116 1272
rect 371016 1232 371022 1244
rect 376110 1232 376116 1244
rect 376168 1232 376174 1284
rect 376478 1232 376484 1284
rect 376536 1272 376542 1284
rect 382366 1272 382372 1284
rect 376536 1244 382372 1272
rect 376536 1232 376542 1244
rect 382366 1232 382372 1244
rect 382424 1232 382430 1284
rect 388622 1232 388628 1284
rect 388680 1272 388686 1284
rect 395338 1272 395344 1284
rect 388680 1244 395344 1272
rect 388680 1232 388686 1244
rect 395338 1232 395344 1244
rect 395396 1232 395402 1284
rect 404078 1232 404084 1284
rect 404136 1272 404142 1284
rect 411898 1272 411904 1284
rect 404136 1244 411904 1272
rect 404136 1232 404142 1244
rect 411898 1232 411904 1244
rect 411956 1232 411962 1284
rect 413922 1232 413928 1284
rect 413980 1272 413986 1284
rect 422570 1272 422576 1284
rect 413980 1244 422576 1272
rect 413980 1232 413986 1244
rect 422570 1232 422576 1244
rect 422628 1232 422634 1284
rect 426158 1232 426164 1284
rect 426216 1272 426222 1284
rect 435174 1272 435180 1284
rect 426216 1244 435180 1272
rect 426216 1232 426222 1244
rect 435174 1232 435180 1244
rect 435232 1232 435238 1284
rect 436002 1232 436008 1284
rect 436060 1272 436066 1284
rect 443840 1272 443868 1312
rect 445846 1300 445852 1312
rect 445904 1300 445910 1352
rect 449342 1300 449348 1352
rect 449400 1340 449406 1352
rect 453206 1340 453212 1352
rect 449400 1312 453212 1340
rect 449400 1300 449406 1312
rect 453206 1300 453212 1312
rect 453264 1300 453270 1352
rect 455690 1340 455696 1352
rect 453408 1312 455696 1340
rect 436060 1244 443868 1272
rect 436060 1232 436066 1244
rect 444926 1232 444932 1284
rect 444984 1272 444990 1284
rect 453408 1272 453436 1312
rect 455690 1300 455696 1312
rect 455748 1300 455754 1352
rect 462590 1300 462596 1352
rect 462648 1340 462654 1352
rect 474182 1340 474188 1352
rect 462648 1312 474188 1340
rect 462648 1300 462654 1312
rect 474182 1300 474188 1312
rect 474240 1300 474246 1352
rect 475838 1300 475844 1352
rect 475896 1340 475902 1352
rect 488810 1340 488816 1352
rect 475896 1312 488816 1340
rect 475896 1300 475902 1312
rect 488810 1300 488816 1312
rect 488868 1300 488874 1352
rect 493502 1300 493508 1352
rect 493560 1340 493566 1352
rect 507302 1340 507308 1352
rect 493560 1312 507308 1340
rect 493560 1300 493566 1312
rect 507302 1300 507308 1312
rect 507360 1300 507366 1352
rect 526622 1300 526628 1352
rect 526680 1340 526686 1352
rect 535546 1340 535552 1352
rect 526680 1312 535552 1340
rect 526680 1300 526686 1312
rect 535546 1300 535552 1312
rect 535604 1300 535610 1352
rect 539870 1300 539876 1352
rect 539928 1340 539934 1352
rect 556982 1340 556988 1352
rect 539928 1312 556988 1340
rect 539928 1300 539934 1312
rect 556982 1300 556988 1312
rect 557040 1300 557046 1352
rect 444984 1244 453436 1272
rect 444984 1232 444990 1244
rect 454862 1232 454868 1284
rect 454920 1272 454926 1284
rect 465994 1272 466000 1284
rect 454920 1244 466000 1272
rect 454920 1232 454926 1244
rect 465994 1232 466000 1244
rect 466052 1232 466058 1284
rect 469122 1232 469128 1284
rect 469180 1272 469186 1284
rect 481358 1272 481364 1284
rect 469180 1244 481364 1272
rect 469180 1232 469186 1244
rect 481358 1232 481364 1244
rect 481416 1232 481422 1284
rect 495710 1232 495716 1284
rect 495768 1272 495774 1284
rect 509694 1272 509700 1284
rect 495768 1244 509700 1272
rect 495768 1232 495774 1244
rect 509694 1232 509700 1244
rect 509752 1232 509758 1284
rect 510062 1232 510068 1284
rect 510120 1272 510126 1284
rect 520182 1272 520188 1284
rect 510120 1244 520188 1272
rect 510120 1232 510126 1244
rect 520182 1232 520188 1244
rect 520240 1232 520246 1284
rect 524322 1232 524328 1284
rect 524380 1272 524386 1284
rect 532602 1272 532608 1284
rect 524380 1244 532608 1272
rect 524380 1232 524386 1244
rect 532602 1232 532608 1244
rect 532660 1232 532666 1284
rect 68830 1164 68836 1216
rect 68888 1204 68894 1216
rect 79410 1204 79416 1216
rect 68888 1176 79416 1204
rect 68888 1164 68894 1176
rect 79410 1164 79416 1176
rect 79468 1164 79474 1216
rect 268838 1164 268844 1216
rect 268896 1204 268902 1216
rect 270402 1204 270408 1216
rect 268896 1176 270408 1204
rect 268896 1164 268902 1176
rect 270402 1164 270408 1176
rect 270460 1164 270466 1216
rect 359918 1164 359924 1216
rect 359976 1204 359982 1216
rect 364610 1204 364616 1216
rect 359976 1176 364616 1204
rect 359976 1164 359982 1176
rect 364610 1164 364616 1176
rect 364668 1164 364674 1216
rect 368750 1164 368756 1216
rect 368808 1204 368814 1216
rect 373902 1204 373908 1216
rect 368808 1176 373908 1204
rect 368808 1164 368814 1176
rect 373902 1164 373908 1176
rect 373960 1164 373966 1216
rect 378686 1164 378692 1216
rect 378744 1204 378750 1216
rect 384390 1204 384396 1216
rect 378744 1176 384396 1204
rect 378744 1164 378750 1176
rect 384390 1164 384396 1176
rect 384448 1164 384454 1216
rect 387518 1164 387524 1216
rect 387576 1204 387582 1216
rect 394234 1204 394240 1216
rect 387576 1176 394240 1204
rect 387576 1164 387582 1176
rect 394234 1164 394240 1176
rect 394292 1164 394298 1216
rect 395246 1164 395252 1216
rect 395304 1204 395310 1216
rect 402514 1204 402520 1216
rect 395304 1176 402520 1204
rect 395304 1164 395310 1176
rect 402514 1164 402520 1176
rect 402572 1164 402578 1216
rect 420638 1164 420644 1216
rect 420696 1204 420702 1216
rect 429286 1204 429292 1216
rect 420696 1176 429292 1204
rect 420696 1164 420702 1176
rect 429286 1164 429292 1176
rect 429344 1164 429350 1216
rect 434990 1164 434996 1216
rect 435048 1204 435054 1216
rect 445018 1204 445024 1216
rect 435048 1176 445024 1204
rect 435048 1164 435054 1176
rect 445018 1164 445024 1176
rect 445076 1164 445082 1216
rect 445956 1176 448652 1204
rect 352190 1096 352196 1148
rect 352248 1136 352254 1148
rect 356330 1136 356336 1148
rect 352248 1108 356336 1136
rect 352248 1096 352254 1108
rect 356330 1096 356336 1108
rect 356388 1096 356394 1148
rect 361022 1096 361028 1148
rect 361080 1136 361086 1148
rect 365438 1136 365444 1148
rect 361080 1108 365444 1136
rect 361080 1096 361086 1108
rect 365438 1096 365444 1108
rect 365496 1096 365502 1148
rect 369762 1096 369768 1148
rect 369820 1136 369826 1148
rect 375282 1136 375288 1148
rect 369820 1108 375288 1136
rect 369820 1096 369826 1108
rect 375282 1096 375288 1108
rect 375340 1096 375346 1148
rect 379790 1096 379796 1148
rect 379848 1136 379854 1148
rect 385954 1136 385960 1148
rect 379848 1108 385960 1136
rect 379848 1096 379854 1108
rect 385954 1096 385960 1108
rect 386012 1096 386018 1148
rect 397362 1096 397368 1148
rect 397420 1136 397426 1148
rect 404814 1136 404820 1148
rect 397420 1108 404820 1136
rect 397420 1096 397426 1108
rect 404814 1096 404820 1108
rect 404872 1096 404878 1148
rect 412910 1096 412916 1148
rect 412968 1136 412974 1148
rect 421374 1136 421380 1148
rect 412968 1108 421380 1136
rect 412968 1096 412974 1108
rect 421374 1096 421380 1108
rect 421432 1096 421438 1148
rect 422846 1096 422852 1148
rect 422904 1136 422910 1148
rect 431862 1136 431868 1148
rect 422904 1108 431868 1136
rect 422904 1096 422910 1108
rect 431862 1096 431868 1108
rect 431920 1096 431926 1148
rect 438302 1096 438308 1148
rect 438360 1136 438366 1148
rect 445754 1136 445760 1148
rect 438360 1108 445760 1136
rect 438360 1096 438366 1108
rect 445754 1096 445760 1108
rect 445812 1096 445818 1148
rect 355502 1028 355508 1080
rect 355560 1068 355566 1080
rect 359918 1068 359924 1080
rect 355560 1040 359924 1068
rect 355560 1028 355566 1040
rect 359918 1028 359924 1040
rect 359976 1028 359982 1080
rect 366542 1028 366548 1080
rect 366600 1068 366606 1080
rect 371326 1068 371332 1080
rect 366600 1040 371332 1068
rect 366600 1028 366606 1040
rect 371326 1028 371332 1040
rect 371384 1028 371390 1080
rect 373166 1028 373172 1080
rect 373224 1068 373230 1080
rect 378502 1068 378508 1080
rect 373224 1040 378508 1068
rect 373224 1028 373230 1040
rect 378502 1028 378508 1040
rect 378560 1028 378566 1080
rect 394142 1028 394148 1080
rect 394200 1068 394206 1080
rect 401318 1068 401324 1080
rect 394200 1040 401324 1068
rect 394200 1028 394206 1040
rect 401318 1028 401324 1040
rect 401376 1028 401382 1080
rect 424962 1028 424968 1080
rect 425020 1068 425026 1080
rect 434070 1068 434076 1080
rect 425020 1040 434076 1068
rect 425020 1028 425026 1040
rect 434070 1028 434076 1040
rect 434128 1028 434134 1080
rect 442718 1028 442724 1080
rect 442776 1068 442782 1080
rect 445956 1068 445984 1176
rect 448624 1136 448652 1176
rect 450446 1164 450452 1216
rect 450504 1204 450510 1216
rect 461578 1204 461584 1216
rect 450504 1176 461584 1204
rect 450504 1164 450510 1176
rect 461578 1164 461584 1176
rect 461636 1164 461642 1216
rect 482462 1164 482468 1216
rect 482520 1204 482526 1216
rect 495526 1204 495532 1216
rect 482520 1176 495532 1204
rect 482520 1164 482526 1176
rect 495526 1164 495532 1176
rect 495584 1164 495590 1216
rect 506750 1164 506756 1216
rect 506808 1204 506814 1216
rect 514846 1204 514852 1216
rect 506808 1176 514852 1204
rect 506808 1164 506814 1176
rect 514846 1164 514852 1176
rect 514904 1164 514910 1216
rect 528830 1164 528836 1216
rect 528888 1204 528894 1216
rect 545482 1204 545488 1216
rect 528888 1176 545488 1204
rect 528888 1164 528894 1176
rect 545482 1164 545488 1176
rect 545540 1164 545546 1216
rect 453298 1136 453304 1148
rect 448624 1108 453304 1136
rect 453298 1096 453304 1108
rect 453356 1096 453362 1148
rect 455966 1096 455972 1148
rect 456024 1136 456030 1148
rect 467466 1136 467472 1148
rect 456024 1108 467472 1136
rect 456024 1096 456030 1108
rect 467466 1096 467472 1108
rect 467524 1096 467530 1148
rect 474642 1096 474648 1148
rect 474700 1136 474706 1148
rect 487246 1136 487252 1148
rect 474700 1108 487252 1136
rect 474700 1096 474706 1108
rect 487246 1096 487252 1108
rect 487304 1096 487310 1148
rect 487982 1096 487988 1148
rect 488040 1136 488046 1148
rect 501414 1136 501420 1148
rect 488040 1108 501420 1136
rect 488040 1096 488046 1108
rect 501414 1096 501420 1108
rect 501472 1096 501478 1148
rect 507762 1096 507768 1148
rect 507820 1136 507826 1148
rect 514754 1136 514760 1148
rect 507820 1108 514760 1136
rect 507820 1096 507826 1108
rect 514754 1096 514760 1108
rect 514812 1096 514818 1148
rect 533246 1096 533252 1148
rect 533304 1136 533310 1148
rect 541526 1136 541532 1148
rect 533304 1108 541532 1136
rect 533304 1096 533310 1108
rect 541526 1096 541532 1108
rect 541584 1096 541590 1148
rect 442776 1040 445984 1068
rect 442776 1028 442782 1040
rect 446030 1028 446036 1080
rect 446088 1068 446094 1080
rect 446088 1040 448652 1068
rect 446088 1028 446094 1040
rect 345566 960 345572 1012
rect 345624 1000 345630 1012
rect 349246 1000 349252 1012
rect 345624 972 349252 1000
rect 345624 960 345630 972
rect 349246 960 349252 972
rect 349304 960 349310 1012
rect 351086 960 351092 1012
rect 351144 1000 351150 1012
rect 355226 1000 355232 1012
rect 351144 972 355232 1000
rect 351144 960 351150 972
rect 355226 960 355232 972
rect 355284 960 355290 1012
rect 362126 960 362132 1012
rect 362184 1000 362190 1012
rect 367002 1000 367008 1012
rect 362184 972 367008 1000
rect 362184 960 362190 972
rect 367002 960 367008 972
rect 367060 960 367066 1012
rect 367646 960 367652 1012
rect 367704 1000 367710 1012
rect 372890 1000 372896 1012
rect 367704 972 372896 1000
rect 367704 960 367710 972
rect 372890 960 372896 972
rect 372948 960 372954 1012
rect 375190 960 375196 1012
rect 375248 1000 375254 1012
rect 381170 1000 381176 1012
rect 375248 972 381176 1000
rect 375248 960 375254 972
rect 381170 960 381176 972
rect 381228 960 381234 1012
rect 419442 960 419448 1012
rect 419500 1000 419506 1012
rect 428458 1000 428464 1012
rect 419500 972 428464 1000
rect 419500 960 419506 972
rect 428458 960 428464 972
rect 428516 960 428522 1012
rect 431678 960 431684 1012
rect 431736 1000 431742 1012
rect 441430 1000 441436 1012
rect 431736 972 441436 1000
rect 431736 960 431742 972
rect 441430 960 441436 972
rect 441488 960 441494 1012
rect 441522 960 441528 1012
rect 441580 1000 441586 1012
rect 448514 1000 448520 1012
rect 441580 972 448520 1000
rect 441580 960 441586 972
rect 448514 960 448520 972
rect 448572 960 448578 1012
rect 19426 892 19432 944
rect 19484 932 19490 944
rect 37458 932 37464 944
rect 19484 904 37464 932
rect 19484 892 19490 904
rect 37458 892 37464 904
rect 37516 892 37522 944
rect 358722 892 358728 944
rect 358780 932 358786 944
rect 363506 932 363512 944
rect 358780 904 363512 932
rect 358780 892 358786 904
rect 363506 892 363512 904
rect 363564 892 363570 944
rect 377582 892 377588 944
rect 377640 932 377646 944
rect 383562 932 383568 944
rect 377640 904 383568 932
rect 377640 892 377646 904
rect 383562 892 383568 904
rect 383620 892 383626 944
rect 416222 892 416228 944
rect 416280 932 416286 944
rect 424962 932 424968 944
rect 416280 904 424968 932
rect 416280 892 416286 904
rect 424962 892 424968 904
rect 425020 892 425026 944
rect 430482 892 430488 944
rect 430540 932 430546 944
rect 430540 904 431954 932
rect 430540 892 430546 904
rect 21818 824 21824 876
rect 21876 864 21882 876
rect 39666 864 39672 876
rect 21876 836 39672 864
rect 21876 824 21882 836
rect 39666 824 39672 836
rect 39724 824 39730 876
rect 337838 824 337844 876
rect 337896 864 337902 876
rect 340966 864 340972 876
rect 337896 836 340972 864
rect 337896 824 337902 836
rect 340966 824 340972 836
rect 341024 824 341030 876
rect 347682 824 347688 876
rect 347740 864 347746 876
rect 351638 864 351644 876
rect 347740 836 351644 864
rect 347740 824 347746 836
rect 351638 824 351644 836
rect 351696 824 351702 876
rect 386322 824 386328 876
rect 386380 864 386386 876
rect 392670 864 392676 876
rect 386380 836 392676 864
rect 386380 824 386386 836
rect 392670 824 392676 836
rect 392728 824 392734 876
rect 421742 824 421748 876
rect 421800 864 421806 876
rect 430850 864 430856 876
rect 421800 836 430856 864
rect 421800 824 421806 836
rect 430850 824 430856 836
rect 430908 824 430914 876
rect 431926 864 431954 904
rect 437198 892 437204 944
rect 437256 932 437262 944
rect 447410 932 447416 944
rect 437256 904 447416 932
rect 437256 892 437262 904
rect 447410 892 447416 904
rect 447468 892 447474 944
rect 448624 932 448652 1040
rect 451550 1028 451556 1080
rect 451608 1068 451614 1080
rect 462406 1068 462412 1080
rect 451608 1040 462412 1068
rect 451608 1028 451614 1040
rect 462406 1028 462412 1040
rect 462464 1028 462470 1080
rect 485682 1028 485688 1080
rect 485740 1068 485746 1080
rect 490098 1068 490104 1080
rect 485740 1040 490104 1068
rect 485740 1028 485746 1040
rect 490098 1028 490104 1040
rect 490156 1028 490162 1080
rect 490190 1028 490196 1080
rect 490248 1068 490254 1080
rect 494790 1068 494796 1080
rect 490248 1040 494796 1068
rect 490248 1028 490254 1040
rect 494790 1028 494796 1040
rect 494848 1028 494854 1080
rect 525518 1028 525524 1080
rect 525576 1068 525582 1080
rect 536834 1068 536840 1080
rect 525576 1040 536840 1068
rect 525576 1028 525582 1040
rect 536834 1028 536840 1040
rect 536892 1028 536898 1080
rect 448698 960 448704 1012
rect 448756 1000 448762 1012
rect 451734 1000 451740 1012
rect 448756 972 451740 1000
rect 448756 960 448762 972
rect 451734 960 451740 972
rect 451792 960 451798 1012
rect 453206 960 453212 1012
rect 453264 1000 453270 1012
rect 453264 972 457024 1000
rect 453264 960 453270 972
rect 456886 932 456892 944
rect 448624 904 456892 932
rect 456886 892 456892 904
rect 456944 892 456950 944
rect 456996 932 457024 972
rect 457070 960 457076 1012
rect 457128 1000 457134 1012
rect 468294 1000 468300 1012
rect 457128 972 468300 1000
rect 457128 960 457134 972
rect 468294 960 468300 972
rect 468352 960 468358 1012
rect 486878 960 486884 1012
rect 486936 1000 486942 1012
rect 500586 1000 500592 1012
rect 486936 972 500592 1000
rect 486936 960 486942 972
rect 500586 960 500592 972
rect 500644 960 500650 1012
rect 501230 960 501236 1012
rect 501288 1000 501294 1012
rect 515490 1000 515496 1012
rect 501288 972 515496 1000
rect 501288 960 501294 972
rect 515490 960 515496 972
rect 515548 960 515554 1012
rect 515582 960 515588 1012
rect 515640 1000 515646 1012
rect 525794 1000 525800 1012
rect 515640 972 525800 1000
rect 515640 960 515646 972
rect 525794 960 525800 972
rect 525852 960 525858 1012
rect 527726 960 527732 1012
rect 527784 1000 527790 1012
rect 544378 1000 544384 1012
rect 527784 972 544384 1000
rect 527784 960 527790 972
rect 544378 960 544384 972
rect 544436 960 544442 1012
rect 460014 932 460020 944
rect 456996 904 460020 932
rect 460014 892 460020 904
rect 460072 892 460078 944
rect 481542 892 481548 944
rect 481600 932 481606 944
rect 481600 904 489914 932
rect 481600 892 481606 904
rect 440326 864 440332 876
rect 431926 836 440332 864
rect 440326 824 440332 836
rect 440384 824 440390 876
rect 447042 824 447048 876
rect 447100 864 447106 876
rect 458082 864 458088 876
rect 447100 836 458088 864
rect 447100 824 447106 836
rect 458082 824 458088 836
rect 458140 824 458146 876
rect 489886 864 489914 904
rect 494606 892 494612 944
rect 494664 932 494670 944
rect 508866 932 508872 944
rect 494664 904 508872 932
rect 494664 892 494670 904
rect 508866 892 508872 904
rect 508924 892 508930 944
rect 519998 892 520004 944
rect 520056 932 520062 944
rect 536098 932 536104 944
rect 520056 904 536104 932
rect 520056 892 520062 904
rect 536098 892 536104 904
rect 536156 892 536162 944
rect 494698 864 494704 876
rect 489886 836 494704 864
rect 494698 824 494704 836
rect 494756 824 494762 876
rect 494790 824 494796 876
rect 494848 864 494854 876
rect 503806 864 503812 876
rect 494848 836 503812 864
rect 494848 824 494854 836
rect 503806 824 503812 836
rect 503864 824 503870 876
rect 523310 824 523316 876
rect 523368 864 523374 876
rect 532234 864 532240 876
rect 523368 836 532240 864
rect 523368 824 523374 836
rect 532234 824 532240 836
rect 532292 824 532298 876
rect 547598 824 547604 876
rect 547656 864 547662 876
rect 565630 864 565636 876
rect 547656 836 565636 864
rect 547656 824 547662 836
rect 565630 824 565636 836
rect 565688 824 565694 876
rect 8754 756 8760 808
rect 8812 796 8818 808
rect 27522 796 27528 808
rect 8812 768 27528 796
rect 8812 756 8818 768
rect 27522 756 27528 768
rect 27580 756 27586 808
rect 251174 756 251180 808
rect 251232 796 251238 808
rect 253842 796 253848 808
rect 251232 768 253848 796
rect 251232 756 251238 768
rect 253842 756 253848 768
rect 253900 756 253906 808
rect 429470 756 429476 808
rect 429528 796 429534 808
rect 439130 796 439136 808
rect 429528 768 439136 796
rect 429528 756 429534 768
rect 439130 756 439136 768
rect 439188 756 439194 808
rect 440510 756 440516 808
rect 440568 796 440574 808
rect 450906 796 450912 808
rect 440568 768 450912 796
rect 440568 756 440574 768
rect 450906 756 450912 768
rect 450964 756 450970 808
rect 483566 756 483572 808
rect 483624 796 483630 808
rect 497090 796 497096 808
rect 483624 768 497096 796
rect 483624 756 483630 768
rect 497090 756 497096 768
rect 497148 756 497154 808
rect 514478 756 514484 808
rect 514536 796 514542 808
rect 529750 796 529756 808
rect 514536 768 529756 796
rect 514536 756 514542 768
rect 529750 756 529756 768
rect 529808 756 529814 808
rect 532142 756 532148 808
rect 532200 796 532206 808
rect 548702 796 548708 808
rect 532200 768 548708 796
rect 532200 756 532206 768
rect 548702 756 548708 768
rect 548760 756 548766 808
rect 550910 756 550916 808
rect 550968 796 550974 808
rect 569126 796 569132 808
rect 550968 768 569132 796
rect 550968 756 550974 768
rect 569126 756 569132 768
rect 569184 756 569190 808
rect 17034 688 17040 740
rect 17092 728 17098 740
rect 35250 728 35256 740
rect 17092 700 35256 728
rect 17092 688 17098 700
rect 35250 688 35256 700
rect 35308 688 35314 740
rect 432782 688 432788 740
rect 432840 728 432846 740
rect 442626 728 442632 740
rect 432840 700 442632 728
rect 432840 688 432846 700
rect 442626 688 442632 700
rect 442684 688 442690 740
rect 443822 688 443828 740
rect 443880 728 443886 740
rect 454126 728 454132 740
rect 443880 700 454132 728
rect 443880 688 443886 700
rect 454126 688 454132 700
rect 454184 688 454190 740
rect 468110 688 468116 740
rect 468168 728 468174 740
rect 480530 728 480536 740
rect 468168 700 480536 728
rect 468168 688 468174 700
rect 480530 688 480536 700
rect 480588 688 480594 740
rect 489086 688 489092 740
rect 489144 728 489150 740
rect 502978 728 502984 740
rect 489144 700 502984 728
rect 489144 688 489150 700
rect 502978 688 502984 700
rect 503036 688 503042 740
rect 522206 688 522212 740
rect 522264 728 522270 740
rect 538214 728 538220 740
rect 522264 700 538220 728
rect 522264 688 522270 700
rect 538214 688 538220 700
rect 538272 688 538278 740
rect 540882 688 540888 740
rect 540940 728 540946 740
rect 558546 728 558552 740
rect 540940 700 558552 728
rect 540940 688 540946 700
rect 558546 688 558552 700
rect 558604 688 558610 740
rect 15930 620 15936 672
rect 15988 660 15994 672
rect 34146 660 34152 672
rect 15988 632 34152 660
rect 15988 620 15994 632
rect 34146 620 34152 632
rect 34204 620 34210 672
rect 35986 620 35992 672
rect 36044 660 36050 672
rect 52914 660 52920 672
rect 36044 632 52920 660
rect 36044 620 36050 632
rect 52914 620 52920 632
rect 52972 620 52978 672
rect 400122 660 400128 672
rect 393286 632 400128 660
rect 11146 552 11152 604
rect 11204 592 11210 604
rect 29730 592 29736 604
rect 11204 564 29736 592
rect 11204 552 11210 564
rect 29730 552 29736 564
rect 29788 552 29794 604
rect 39574 552 39580 604
rect 39632 592 39638 604
rect 56226 592 56232 604
rect 39632 564 56232 592
rect 39632 552 39638 564
rect 56226 552 56232 564
rect 56284 552 56290 604
rect 384206 552 384212 604
rect 384264 592 384270 604
rect 390646 592 390652 604
rect 384264 564 390652 592
rect 384264 552 384270 564
rect 390646 552 390652 564
rect 390704 552 390710 604
rect 393038 552 393044 604
rect 393096 592 393102 604
rect 393286 592 393314 632
rect 400122 620 400128 632
rect 400180 620 400186 672
rect 401870 620 401876 672
rect 401928 660 401934 672
rect 409230 660 409236 672
rect 401928 632 409236 660
rect 401928 620 401934 632
rect 409230 620 409236 632
rect 409288 620 409294 672
rect 417878 660 417884 672
rect 412606 632 417884 660
rect 393096 564 393314 592
rect 393096 552 393102 564
rect 397730 552 397736 604
rect 397788 552 397794 604
rect 408402 552 408408 604
rect 408460 552 408466 604
rect 409598 552 409604 604
rect 409656 592 409662 604
rect 412606 592 412634 632
rect 417878 620 417884 632
rect 417936 620 417942 672
rect 427262 620 427268 672
rect 427320 660 427326 672
rect 436738 660 436744 672
rect 427320 632 436744 660
rect 427320 620 427326 632
rect 436738 620 436744 632
rect 436796 620 436802 672
rect 448238 620 448244 672
rect 448296 660 448302 672
rect 459186 660 459192 672
rect 448296 632 459192 660
rect 448296 620 448302 632
rect 459186 620 459192 632
rect 459244 620 459250 672
rect 459278 620 459284 672
rect 459336 660 459342 672
rect 471054 660 471060 672
rect 459336 632 471060 660
rect 459336 620 459342 632
rect 471054 620 471060 632
rect 471112 620 471118 672
rect 471422 620 471428 672
rect 471480 660 471486 672
rect 479518 660 479524 672
rect 471480 632 479524 660
rect 471480 620 471486 632
rect 479518 620 479524 632
rect 479576 620 479582 672
rect 480162 620 480168 672
rect 480220 660 480226 672
rect 493134 660 493140 672
rect 480220 632 493140 660
rect 480220 620 480226 632
rect 493134 620 493140 632
rect 493192 620 493198 672
rect 502242 620 502248 672
rect 502300 660 502306 672
rect 517146 660 517152 672
rect 502300 632 517152 660
rect 502300 620 502306 632
rect 517146 620 517152 632
rect 517204 620 517210 672
rect 542078 620 542084 672
rect 542136 660 542142 672
rect 559742 660 559748 672
rect 542136 632 559748 660
rect 542136 620 542142 632
rect 559742 620 559748 632
rect 559800 620 559806 672
rect 563238 660 563244 672
rect 561968 632 563244 660
rect 409656 564 412634 592
rect 409656 552 409662 564
rect 416682 552 416688 604
rect 416740 552 416746 604
rect 433886 552 433892 604
rect 433944 592 433950 604
rect 443454 592 443460 604
rect 433944 564 443460 592
rect 433944 552 433950 564
rect 443454 552 443460 564
rect 443512 552 443518 604
rect 443730 552 443736 604
rect 443788 592 443794 604
rect 449802 592 449808 604
rect 443788 564 449808 592
rect 443788 552 443794 564
rect 449802 552 449808 564
rect 449860 552 449866 604
rect 461486 552 461492 604
rect 461544 592 461550 604
rect 473446 592 473452 604
rect 461544 564 473452 592
rect 461544 552 461550 564
rect 473446 552 473452 564
rect 473504 552 473510 604
rect 491202 552 491208 604
rect 491260 592 491266 604
rect 505370 592 505376 604
rect 491260 564 505376 592
rect 491260 552 491266 564
rect 505370 552 505376 564
rect 505428 552 505434 604
rect 508958 552 508964 604
rect 509016 592 509022 604
rect 524230 592 524236 604
rect 509016 564 524236 592
rect 509016 552 509022 564
rect 524230 552 524236 564
rect 524288 552 524294 604
rect 545390 552 545396 604
rect 545448 592 545454 604
rect 561968 592 561996 632
rect 563238 620 563244 632
rect 563296 620 563302 672
rect 545448 564 561996 592
rect 545448 552 545454 564
rect 562042 552 562048 604
rect 562100 552 562106 604
rect 18046 484 18052 536
rect 18104 524 18110 536
rect 36354 524 36360 536
rect 18104 496 36360 524
rect 18104 484 18110 496
rect 36354 484 36360 496
rect 36412 484 36418 536
rect 38562 484 38568 536
rect 38620 524 38626 536
rect 55122 524 55128 536
rect 38620 496 55128 524
rect 38620 484 38626 496
rect 55122 484 55128 496
rect 55180 484 55186 536
rect 390830 484 390836 536
rect 390888 524 390894 536
rect 397748 524 397776 552
rect 390888 496 397776 524
rect 390888 484 390894 496
rect 14550 416 14556 468
rect 14608 456 14614 468
rect 33042 456 33048 468
rect 14608 428 33048 456
rect 14608 416 14614 428
rect 33042 416 33048 428
rect 33100 416 33106 468
rect 34606 416 34612 468
rect 34664 456 34670 468
rect 51810 456 51816 468
rect 34664 428 51816 456
rect 34664 416 34670 428
rect 51810 416 51816 428
rect 51868 416 51874 468
rect 381998 416 382004 468
rect 382056 456 382062 468
rect 387886 456 387892 468
rect 382056 428 387892 456
rect 382056 416 382062 428
rect 387886 416 387892 428
rect 387944 416 387950 468
rect 408420 456 408448 552
rect 416700 456 416728 552
rect 470318 484 470324 536
rect 470376 524 470382 536
rect 482462 524 482468 536
rect 470376 496 482468 524
rect 470376 484 470382 496
rect 482462 484 482468 496
rect 482520 484 482526 536
rect 490098 484 490104 536
rect 490156 524 490162 536
rect 499114 524 499120 536
rect 490156 496 499120 524
rect 490156 484 490162 496
rect 499114 484 499120 496
rect 499172 484 499178 536
rect 503438 484 503444 536
rect 503496 524 503502 536
rect 517974 524 517980 536
rect 503496 496 517980 524
rect 503496 484 503502 496
rect 517974 484 517980 496
rect 518032 484 518038 536
rect 544562 484 544568 536
rect 544620 524 544626 536
rect 562060 524 562088 552
rect 544620 496 562088 524
rect 544620 484 544626 496
rect 408420 428 416728 456
rect 464798 416 464804 468
rect 464856 456 464862 468
rect 476574 456 476580 468
rect 464856 428 476580 456
rect 464856 416 464862 428
rect 476574 416 476580 428
rect 476632 416 476638 468
rect 478322 416 478328 468
rect 478380 456 478386 468
rect 490742 456 490748 468
rect 478380 428 490748 456
rect 478380 416 478386 428
rect 490742 416 490748 428
rect 490800 416 490806 468
rect 497918 416 497924 468
rect 497976 456 497982 468
rect 512086 456 512092 468
rect 497976 428 512092 456
rect 497976 416 497982 428
rect 512086 416 512092 428
rect 512144 416 512150 468
rect 516686 416 516692 468
rect 516744 456 516750 468
rect 532142 456 532148 468
rect 516744 428 532148 456
rect 516744 416 516750 428
rect 532142 416 532148 428
rect 532200 416 532206 468
rect 548886 416 548892 468
rect 548944 456 548950 468
rect 567010 456 567016 468
rect 548944 428 567016 456
rect 548944 416 548950 428
rect 567010 416 567016 428
rect 567068 416 567074 468
rect 9766 348 9772 400
rect 9824 388 9830 400
rect 28626 388 28632 400
rect 9824 360 28632 388
rect 9824 348 9830 360
rect 28626 348 28632 360
rect 28684 348 28690 400
rect 32214 348 32220 400
rect 32272 388 32278 400
rect 49602 388 49608 400
rect 32272 360 49608 388
rect 32272 348 32278 360
rect 49602 348 49608 360
rect 49660 348 49666 400
rect 405182 348 405188 400
rect 405240 388 405246 400
rect 412818 388 412824 400
rect 405240 360 412824 388
rect 405240 348 405246 360
rect 412818 348 412824 360
rect 412876 348 412882 400
rect 418430 348 418436 400
rect 418488 388 418494 400
rect 426894 388 426900 400
rect 418488 360 426900 388
rect 418488 348 418494 360
rect 426894 348 426900 360
rect 426952 348 426958 400
rect 453758 348 453764 400
rect 453816 388 453822 400
rect 464982 388 464988 400
rect 453816 360 464988 388
rect 453816 348 453822 360
rect 464982 348 464988 360
rect 465040 348 465046 400
rect 472526 348 472532 400
rect 472584 388 472590 400
rect 472584 360 479288 388
rect 472584 348 472590 360
rect 3234 280 3240 332
rect 3292 320 3298 332
rect 22002 320 22008 332
rect 3292 292 22008 320
rect 3292 280 3298 292
rect 22002 280 22008 292
rect 22060 280 22066 332
rect 22830 280 22836 332
rect 22888 320 22894 332
rect 40494 320 40500 332
rect 22888 292 40500 320
rect 22888 280 22894 292
rect 40494 280 40500 292
rect 40552 280 40558 332
rect 42886 280 42892 332
rect 42944 320 42950 332
rect 59354 320 59360 332
rect 42944 292 59360 320
rect 42944 280 42950 292
rect 59354 280 59360 292
rect 59412 280 59418 332
rect 391658 280 391664 332
rect 391716 320 391722 332
rect 398742 320 398748 332
rect 391716 292 398748 320
rect 391716 280 391722 292
rect 398742 280 398748 292
rect 398800 280 398806 332
rect 400766 280 400772 332
rect 400824 320 400830 332
rect 408586 320 408592 332
rect 400824 292 408592 320
rect 400824 280 400830 292
rect 408586 280 408592 292
rect 408644 280 408650 332
rect 412082 280 412088 332
rect 412140 320 412146 332
rect 420362 320 420368 332
rect 412140 292 420368 320
rect 412140 280 412146 292
rect 420362 280 420368 292
rect 420420 280 420426 332
rect 457898 280 457904 332
rect 457956 320 457962 332
rect 470042 320 470048 332
rect 457956 292 470048 320
rect 457956 280 457962 292
rect 470042 280 470048 292
rect 470100 280 470106 332
rect 479150 280 479156 332
rect 479208 280 479214 332
rect 479260 320 479288 360
rect 479518 348 479524 400
rect 479576 388 479582 400
rect 484210 388 484216 400
rect 479576 360 484216 388
rect 479576 348 479582 360
rect 484210 348 484216 360
rect 484268 348 484274 400
rect 499022 348 499028 400
rect 499080 388 499086 400
rect 513374 388 513380 400
rect 499080 360 513380 388
rect 499080 348 499086 360
rect 513374 348 513380 360
rect 513432 348 513438 400
rect 517790 348 517796 400
rect 517848 388 517854 400
rect 533890 388 533896 400
rect 517848 360 533896 388
rect 517848 348 517854 360
rect 533890 348 533896 360
rect 533948 348 533954 400
rect 534350 348 534356 400
rect 534408 388 534414 400
rect 551094 388 551100 400
rect 534408 360 551100 388
rect 534408 348 534414 360
rect 551094 348 551100 360
rect 551152 348 551158 400
rect 555326 348 555332 400
rect 555384 388 555390 400
rect 573542 388 573548 400
rect 555384 360 573548 388
rect 555384 348 555390 360
rect 573542 348 573548 360
rect 573600 348 573606 400
rect 484854 320 484860 332
rect 479260 292 484860 320
rect 484854 280 484860 292
rect 484912 280 484918 332
rect 504542 280 504548 332
rect 504600 320 504606 332
rect 519722 320 519728 332
rect 504600 292 519728 320
rect 504600 280 504606 292
rect 519722 280 519728 292
rect 519780 280 519786 332
rect 521102 280 521108 332
rect 521160 320 521166 332
rect 537386 320 537392 332
rect 521160 292 537392 320
rect 521160 280 521166 292
rect 537386 280 537392 292
rect 537444 280 537450 332
rect 538766 280 538772 332
rect 538824 320 538830 332
rect 556338 320 556344 332
rect 538824 292 556344 320
rect 538824 280 538830 292
rect 556338 280 556344 292
rect 556396 280 556402 332
rect 557166 280 557172 332
rect 557224 320 557230 332
rect 575934 320 575940 332
rect 557224 292 575940 320
rect 557224 280 557230 292
rect 575934 280 575940 292
rect 575992 280 575998 332
rect 3878 212 3884 264
rect 3936 252 3942 264
rect 23198 252 23204 264
rect 3936 224 23204 252
rect 3936 212 3942 224
rect 23198 212 23204 224
rect 23256 212 23262 264
rect 24578 212 24584 264
rect 24636 252 24642 264
rect 41598 252 41604 264
rect 24636 224 41604 252
rect 24636 212 24642 224
rect 41598 212 41604 224
rect 41656 212 41662 264
rect 42242 212 42248 264
rect 42300 252 42306 264
rect 58158 252 58164 264
rect 42300 224 58164 252
rect 42300 212 42306 224
rect 58158 212 58164 224
rect 58216 212 58222 264
rect 380802 212 380808 264
rect 380860 252 380866 264
rect 386782 252 386788 264
rect 380860 224 386788 252
rect 380860 212 380866 224
rect 386782 212 386788 224
rect 386840 212 386846 264
rect 398558 212 398564 264
rect 398616 252 398622 264
rect 406194 252 406200 264
rect 398616 224 406200 252
rect 398616 212 398622 224
rect 406194 212 406200 224
rect 406252 212 406258 264
rect 410978 212 410984 264
rect 411036 252 411042 264
rect 418614 252 418620 264
rect 411036 224 418620 252
rect 411036 212 411042 224
rect 418614 212 418620 224
rect 418672 212 418678 264
rect 445754 212 445760 264
rect 445812 252 445818 264
rect 448238 252 448244 264
rect 445812 224 448244 252
rect 445812 212 445818 224
rect 448238 212 448244 224
rect 448296 212 448302 264
rect 465902 212 465908 264
rect 465960 252 465966 264
rect 478322 252 478328 264
rect 465960 224 478328 252
rect 465960 212 465966 224
rect 478322 212 478328 224
rect 478380 212 478386 264
rect 479168 252 479196 280
rect 492490 252 492496 264
rect 479168 224 492496 252
rect 492490 212 492496 224
rect 492548 212 492554 264
rect 492582 212 492588 264
rect 492640 252 492646 264
rect 506658 252 506664 264
rect 492640 224 506664 252
rect 492640 212 492646 224
rect 506658 212 506664 224
rect 506716 212 506722 264
rect 511442 212 511448 264
rect 511500 252 511506 264
rect 526254 252 526260 264
rect 511500 224 526260 252
rect 511500 212 511506 224
rect 526254 212 526260 224
rect 526312 212 526318 264
rect 535362 212 535368 264
rect 535420 252 535426 264
rect 552842 252 552848 264
rect 535420 224 552848 252
rect 535420 212 535426 224
rect 552842 212 552848 224
rect 552900 212 552906 264
rect 554222 212 554228 264
rect 554280 252 554286 264
rect 572898 252 572904 264
rect 554280 224 572904 252
rect 554280 212 554286 224
rect 572898 212 572904 224
rect 572956 212 572962 264
rect 8018 144 8024 196
rect 8076 184 8082 196
rect 26326 184 26332 196
rect 8076 156 26332 184
rect 8076 144 8082 156
rect 26326 144 26332 156
rect 26384 144 26390 196
rect 30282 144 30288 196
rect 30340 184 30346 196
rect 47394 184 47400 196
rect 30340 156 47400 184
rect 30340 144 30346 156
rect 47394 144 47400 156
rect 47452 144 47458 196
rect 389726 144 389732 196
rect 389784 184 389790 196
rect 396166 184 396172 196
rect 389784 156 396172 184
rect 389784 144 389790 156
rect 396166 144 396172 156
rect 396224 144 396230 196
rect 399662 144 399668 196
rect 399720 184 399726 196
rect 407022 184 407028 196
rect 399720 156 407028 184
rect 399720 144 399726 156
rect 407022 144 407028 156
rect 407080 144 407086 196
rect 407390 144 407396 196
rect 407448 184 407454 196
rect 415302 184 415308 196
rect 407448 156 415308 184
rect 407448 144 407454 156
rect 415302 144 415308 156
rect 415360 144 415366 196
rect 417326 144 417332 196
rect 417384 184 417390 196
rect 425790 184 425796 196
rect 417384 156 425796 184
rect 417384 144 417390 156
rect 425790 144 425796 156
rect 425848 144 425854 196
rect 452562 144 452568 196
rect 452620 184 452626 196
rect 464154 184 464160 196
rect 452620 156 464160 184
rect 452620 144 452626 156
rect 464154 144 464160 156
rect 464212 144 464218 196
rect 467006 144 467012 196
rect 467064 184 467070 196
rect 478966 184 478972 196
rect 467064 156 478972 184
rect 467064 144 467070 156
rect 478966 144 478972 156
rect 479024 144 479030 196
rect 484670 144 484676 196
rect 484728 184 484734 196
rect 498378 184 498384 196
rect 484728 156 498384 184
rect 484728 144 484734 156
rect 498378 144 498384 156
rect 498436 144 498442 196
rect 505646 144 505652 196
rect 505704 184 505710 196
rect 520366 184 520372 196
rect 505704 156 520372 184
rect 505704 144 505710 156
rect 520366 144 520372 156
rect 520424 144 520430 196
rect 537662 144 537668 196
rect 537720 184 537726 196
rect 554774 184 554780 196
rect 537720 156 554780 184
rect 537720 144 537726 156
rect 554774 144 554780 156
rect 554832 144 554838 196
rect 558822 144 558828 196
rect 558880 184 558886 196
rect 577130 184 577136 196
rect 558880 156 577136 184
rect 558880 144 558886 156
rect 577130 144 577136 156
rect 577188 144 577194 196
rect 1486 76 1492 128
rect 1544 116 1550 128
rect 20898 116 20904 128
rect 1544 88 20904 116
rect 1544 76 1550 88
rect 20898 76 20904 88
rect 20956 76 20962 128
rect 31110 76 31116 128
rect 31168 116 31174 128
rect 48498 116 48504 128
rect 31168 88 48504 116
rect 31168 76 31174 88
rect 48498 76 48504 88
rect 48556 76 48562 128
rect 53558 76 53564 128
rect 53616 116 53622 128
rect 69474 116 69480 128
rect 53616 88 69480 116
rect 53616 76 53622 88
rect 69474 76 69480 88
rect 69532 76 69538 128
rect 354398 76 354404 128
rect 354456 116 354462 128
rect 358906 116 358912 128
rect 354456 88 358912 116
rect 354456 76 354462 88
rect 358906 76 358912 88
rect 358964 76 358970 128
rect 363230 76 363236 128
rect 363288 116 363294 128
rect 367830 116 367836 128
rect 363288 88 367836 116
rect 363288 76 363294 88
rect 367830 76 367836 88
rect 367888 76 367894 128
rect 402882 76 402888 128
rect 402940 116 402946 128
rect 410978 116 410984 128
rect 402940 88 410984 116
rect 402940 76 402946 88
rect 410978 76 410984 88
rect 411036 76 411042 128
rect 460658 76 460664 128
rect 460716 116 460722 128
rect 472434 116 472440 128
rect 460716 88 472440 116
rect 460716 76 460722 88
rect 472434 76 472440 88
rect 472492 76 472498 128
rect 473630 76 473636 128
rect 473688 116 473694 128
rect 486602 116 486608 128
rect 473688 88 486608 116
rect 473688 76 473694 88
rect 486602 76 486608 88
rect 486660 76 486666 128
rect 500126 76 500132 128
rect 500184 116 500190 128
rect 514938 116 514944 128
rect 500184 88 514944 116
rect 500184 76 500190 88
rect 514938 76 514944 88
rect 514996 76 515002 128
rect 518802 76 518808 128
rect 518860 116 518866 128
rect 534534 116 534540 128
rect 518860 88 534540 116
rect 518860 76 518866 88
rect 534534 76 534540 88
rect 534592 76 534598 128
rect 546402 76 546408 128
rect 546460 116 546466 128
rect 564618 116 564624 128
rect 546460 88 564624 116
rect 546460 76 546466 88
rect 564618 76 564624 88
rect 564676 76 564682 128
rect 382 8 388 60
rect 440 48 446 60
rect 19794 48 19800 60
rect 440 20 19800 48
rect 440 8 446 20
rect 19794 8 19800 20
rect 19852 8 19858 60
rect 20438 8 20444 60
rect 20496 48 20502 60
rect 38194 48 38200 60
rect 20496 20 38200 48
rect 20496 8 20502 20
rect 38194 8 38200 20
rect 38252 8 38258 60
rect 45278 8 45284 60
rect 45336 48 45342 60
rect 61746 48 61752 60
rect 45336 20 61752 48
rect 45336 8 45342 20
rect 61746 8 61752 20
rect 61804 8 61810 60
rect 344738 8 344744 60
rect 344796 48 344802 60
rect 348234 48 348240 60
rect 344796 20 348240 48
rect 344796 8 344802 20
rect 348234 8 348240 20
rect 348292 8 348298 60
rect 383102 8 383108 60
rect 383160 48 383166 60
rect 389634 48 389640 60
rect 383160 20 389640 48
rect 383160 8 383166 20
rect 389634 8 389640 20
rect 389692 8 389698 60
rect 423950 8 423956 60
rect 424008 48 424014 60
rect 433426 48 433432 60
rect 424008 20 433432 48
rect 424008 8 424014 20
rect 433426 8 433432 20
rect 433484 8 433490 60
rect 463602 8 463608 60
rect 463660 48 463666 60
rect 475930 48 475936 60
rect 463660 20 475936 48
rect 463660 8 463666 20
rect 475930 8 475936 20
rect 475988 8 475994 60
rect 477218 8 477224 60
rect 477276 48 477282 60
rect 490098 48 490104 60
rect 477276 20 490104 48
rect 477276 8 477282 20
rect 490098 8 490104 20
rect 490156 8 490162 60
rect 496722 8 496728 60
rect 496780 48 496786 60
rect 511442 48 511448 60
rect 496780 20 511448 48
rect 496780 8 496786 20
rect 511442 8 511448 20
rect 511500 8 511506 60
rect 512638 8 512644 60
rect 512696 48 512702 60
rect 528002 48 528008 60
rect 512696 20 528008 48
rect 512696 8 512702 20
rect 528002 8 528008 20
rect 528060 8 528066 60
rect 531038 8 531044 60
rect 531096 48 531102 60
rect 548058 48 548064 60
rect 531096 20 548064 48
rect 531096 8 531102 20
rect 548058 8 548064 20
rect 548116 8 548122 60
rect 551922 8 551928 60
rect 551980 48 551986 60
rect 570506 48 570512 60
rect 551980 20 570512 48
rect 551980 8 551986 20
rect 570506 8 570512 20
rect 570564 8 570570 60
<< via1 >>
rect 186504 702992 186556 703044
rect 188436 702992 188488 703044
rect 235172 702992 235224 703044
rect 236184 702992 236236 703044
rect 522764 702992 522816 703044
rect 527088 702992 527140 703044
rect 570512 702992 570564 703044
rect 575848 702992 575900 703044
rect 490932 702720 490984 702772
rect 494796 702720 494848 702772
rect 538680 702720 538732 702772
rect 543464 702720 543516 702772
rect 24308 702448 24360 702500
rect 29276 702448 29328 702500
rect 218980 702448 219032 702500
rect 220268 702448 220320 702500
rect 459100 702448 459152 702500
rect 462320 702448 462372 702500
rect 506848 702448 506900 702500
rect 510988 702448 511040 702500
rect 554596 702448 554648 702500
rect 559656 702448 559708 702500
rect 8116 700952 8168 701004
rect 13084 700952 13136 701004
rect 40500 700952 40552 701004
rect 44916 700952 44968 701004
rect 56784 700952 56836 701004
rect 60740 700952 60792 701004
rect 72976 700952 73028 701004
rect 76748 700952 76800 701004
rect 89168 700952 89220 701004
rect 92572 700952 92624 701004
rect 105452 700952 105504 701004
rect 108580 700952 108632 701004
rect 121644 700952 121696 701004
rect 124404 700952 124456 701004
rect 137836 700952 137888 701004
rect 140412 700952 140464 701004
rect 154120 700952 154172 701004
rect 156236 700952 156288 701004
rect 170312 700952 170364 701004
rect 172428 700952 172480 701004
rect 202788 700952 202840 701004
rect 204260 700952 204312 701004
rect 348056 700952 348108 701004
rect 348792 700952 348844 701004
rect 363880 700952 363932 701004
rect 364984 700952 365036 701004
rect 379336 700952 379388 701004
rect 381176 700952 381228 701004
rect 395712 700952 395764 701004
rect 397460 700952 397512 701004
rect 411720 700952 411772 701004
rect 413652 700952 413704 701004
rect 427544 700952 427596 701004
rect 429844 700952 429896 701004
rect 443552 700952 443604 701004
rect 446128 700952 446180 701004
rect 475384 700952 475436 701004
rect 478512 700952 478564 701004
rect 65524 3816 65576 3868
rect 80244 3816 80296 3868
rect 97632 3816 97684 3868
rect 101220 3816 101272 3868
rect 56048 3748 56100 3800
rect 71412 3748 71464 3800
rect 90088 3748 90140 3800
rect 103428 3748 103480 3800
rect 104348 3748 104400 3800
rect 52552 3680 52604 3732
rect 68100 3680 68152 3732
rect 71872 3680 71924 3732
rect 85764 3680 85816 3732
rect 86868 3680 86920 3732
rect 100116 3680 100168 3732
rect 106648 3680 106700 3732
rect 48964 3612 49016 3664
rect 64788 3612 64840 3664
rect 66720 3612 66772 3664
rect 81440 3612 81492 3664
rect 84476 3612 84528 3664
rect 97908 3612 97960 3664
rect 60832 3544 60884 3596
rect 75920 3544 75972 3596
rect 76288 3544 76340 3596
rect 90180 3544 90232 3596
rect 54944 3476 54996 3528
rect 70308 3476 70360 3528
rect 71504 3476 71556 3528
rect 71872 3476 71924 3528
rect 72976 3476 73028 3528
rect 86960 3476 87012 3528
rect 87788 3476 87840 3528
rect 97632 3544 97684 3596
rect 97448 3476 97500 3528
rect 110052 3612 110104 3664
rect 116676 3680 116728 3732
rect 118884 3612 118936 3664
rect 125968 3612 126020 3664
rect 136548 3612 136600 3664
rect 143632 3612 143684 3664
rect 153200 3612 153252 3664
rect 108488 3544 108540 3596
rect 119988 3544 120040 3596
rect 122288 3544 122340 3596
rect 133236 3544 133288 3596
rect 142528 3544 142580 3596
rect 152004 3544 152056 3596
rect 98644 3476 98696 3528
rect 51356 3408 51408 3460
rect 66996 3408 67048 3460
rect 70124 3408 70176 3460
rect 84660 3408 84712 3460
rect 89536 3408 89588 3460
rect 102324 3408 102376 3460
rect 110512 3476 110564 3528
rect 122380 3476 122432 3528
rect 129372 3476 129424 3528
rect 139860 3476 139912 3528
rect 141608 3476 141660 3528
rect 150900 3476 150952 3528
rect 111156 3408 111208 3460
rect 117596 3408 117648 3460
rect 128820 3408 128872 3460
rect 63224 3340 63276 3392
rect 78036 3340 78088 3392
rect 83280 3340 83332 3392
rect 92940 3340 92992 3392
rect 93952 3340 94004 3392
rect 62028 3272 62080 3324
rect 76932 3272 76984 3324
rect 82084 3272 82136 3324
rect 95700 3272 95752 3324
rect 58808 3204 58860 3256
rect 73620 3204 73672 3256
rect 77392 3204 77444 3256
rect 91284 3204 91336 3256
rect 96252 3204 96304 3256
rect 101036 3340 101088 3392
rect 113364 3340 113416 3392
rect 116400 3340 116452 3392
rect 121552 3340 121604 3392
rect 128176 3340 128228 3392
rect 138756 3408 138808 3460
rect 130568 3340 130620 3392
rect 140688 3340 140740 3392
rect 103336 3272 103388 3324
rect 115572 3272 115624 3324
rect 119896 3272 119948 3324
rect 131028 3272 131080 3324
rect 140044 3272 140096 3324
rect 149796 3408 149848 3460
rect 56968 3136 57020 3188
rect 72516 3136 72568 3188
rect 73804 3136 73856 3188
rect 87972 3136 88024 3188
rect 92848 3136 92900 3188
rect 106740 3204 106792 3256
rect 111616 3204 111668 3256
rect 123300 3204 123352 3256
rect 123760 3204 123812 3256
rect 134340 3204 134392 3256
rect 137652 3204 137704 3256
rect 147588 3340 147640 3392
rect 154028 3340 154080 3392
rect 163044 3340 163096 3392
rect 166080 3340 166132 3392
rect 174084 3340 174136 3392
rect 183744 3340 183796 3392
rect 190644 3340 190696 3392
rect 553308 3340 553360 3392
rect 571524 3340 571576 3392
rect 145932 3272 145984 3324
rect 155316 3272 155368 3324
rect 155776 3272 155828 3324
rect 164240 3272 164292 3324
rect 164884 3272 164936 3324
rect 172980 3272 173032 3324
rect 176752 3272 176804 3324
rect 184020 3272 184072 3324
rect 184940 3272 184992 3324
rect 151820 3204 151872 3256
rect 160836 3204 160888 3256
rect 162492 3204 162544 3256
rect 170772 3204 170824 3256
rect 40960 3068 41012 3120
rect 57060 3068 57112 3120
rect 80888 3068 80940 3120
rect 94596 3068 94648 3120
rect 108948 3136 109000 3188
rect 109408 3136 109460 3188
rect 121092 3136 121144 3188
rect 132132 3136 132184 3188
rect 136456 3136 136508 3188
rect 146208 3136 146260 3188
rect 105636 3068 105688 3120
rect 106096 3068 106148 3120
rect 117780 3068 117832 3120
rect 121184 3068 121236 3120
rect 121552 3068 121604 3120
rect 127716 3068 127768 3120
rect 131764 3068 131816 3120
rect 142068 3068 142120 3120
rect 144736 3068 144788 3120
rect 154212 3136 154264 3188
rect 156328 3136 156380 3188
rect 165252 3136 165304 3188
rect 165712 3136 165764 3188
rect 171876 3204 171928 3256
rect 173164 3204 173216 3256
rect 180892 3204 180944 3256
rect 181444 3204 181496 3256
rect 188436 3204 188488 3256
rect 550088 3272 550140 3324
rect 568028 3272 568080 3324
rect 191840 3204 191892 3256
rect 174268 3136 174320 3188
rect 149520 3068 149572 3120
rect 158720 3068 158772 3120
rect 160192 3068 160244 3120
rect 168564 3068 168616 3120
rect 50160 3000 50212 3052
rect 65892 3000 65944 3052
rect 69112 3000 69164 3052
rect 83556 3000 83608 3052
rect 26608 2932 26660 2984
rect 44088 2932 44140 2984
rect 44272 2932 44324 2984
rect 27712 2864 27764 2916
rect 45192 2864 45244 2916
rect 47860 2932 47912 2984
rect 63408 2932 63460 2984
rect 67916 2932 67968 2984
rect 77116 2932 77168 2984
rect 78588 2932 78640 2984
rect 92388 3000 92440 3052
rect 60648 2864 60700 2916
rect 33600 2796 33652 2848
rect 50712 2796 50764 2848
rect 59636 2796 59688 2848
rect 75000 2864 75052 2916
rect 75368 2864 75420 2916
rect 85488 2864 85540 2916
rect 64328 2796 64380 2848
rect 68836 2796 68888 2848
rect 79692 2796 79744 2848
rect 88984 2932 89036 2984
rect 85672 2864 85724 2916
rect 95148 3000 95200 3052
rect 104532 3000 104584 3052
rect 112812 3000 112864 3052
rect 124404 3000 124456 3052
rect 125048 3000 125100 3052
rect 135168 3000 135220 3052
rect 135904 3000 135956 3052
rect 145380 3000 145432 3052
rect 147128 3000 147180 3052
rect 156420 3000 156472 3052
rect 159272 3000 159324 3052
rect 167460 3000 167512 3052
rect 168380 3000 168432 3052
rect 176292 3068 176344 3120
rect 179052 3136 179104 3188
rect 186320 3136 186372 3188
rect 190828 3136 190880 3188
rect 197360 3204 197412 3256
rect 214472 3204 214524 3256
rect 219348 3204 219400 3256
rect 530032 3204 530084 3256
rect 546684 3204 546736 3256
rect 556712 3204 556764 3256
rect 575112 3204 575164 3256
rect 196808 3136 196860 3188
rect 202880 3136 202932 3188
rect 209872 3136 209924 3188
rect 214932 3136 214984 3188
rect 220452 3136 220504 3188
rect 224868 3136 224920 3188
rect 561128 3136 561180 3188
rect 579804 3136 579856 3188
rect 181812 3068 181864 3120
rect 186136 3068 186188 3120
rect 192852 3068 192904 3120
rect 193312 3068 193364 3120
rect 199476 3068 199528 3120
rect 200304 3068 200356 3120
rect 206100 3068 206152 3120
rect 206192 3068 206244 3120
rect 211620 3068 211672 3120
rect 216864 3068 216916 3120
rect 221556 3068 221608 3120
rect 231032 3068 231084 3120
rect 234804 3068 234856 3120
rect 239312 3068 239364 3120
rect 242532 3068 242584 3120
rect 532608 3068 532660 3120
rect 540796 3068 540848 3120
rect 563152 3068 563204 3120
rect 582196 3068 582248 3120
rect 91928 2796 91980 2848
rect 102232 2932 102284 2984
rect 95056 2864 95108 2916
rect 107844 2864 107896 2916
rect 114008 2932 114060 2984
rect 125600 2932 125652 2984
rect 134156 2932 134208 2984
rect 144552 2932 144604 2984
rect 114560 2864 114612 2916
rect 115204 2864 115256 2916
rect 126612 2864 126664 2916
rect 126980 2864 127032 2916
rect 137928 2864 137980 2916
rect 138848 2864 138900 2916
rect 148968 2932 149020 2984
rect 153016 2932 153068 2984
rect 162216 2932 162268 2984
rect 163688 2932 163740 2984
rect 165712 2932 165764 2984
rect 167184 2932 167236 2984
rect 175280 3000 175332 3052
rect 175832 3000 175884 3052
rect 182916 3000 182968 3052
rect 188528 3000 188580 3052
rect 195060 3000 195112 3052
rect 195612 3000 195664 3052
rect 201684 3000 201736 3052
rect 171968 2932 172020 2984
rect 179880 2932 179932 2984
rect 182548 2932 182600 2984
rect 189540 2932 189592 2984
rect 189724 2932 189776 2984
rect 196440 2932 196492 2984
rect 201500 2932 201552 2984
rect 206928 3000 206980 3052
rect 210976 3000 211028 3052
rect 216036 3000 216088 3052
rect 218060 3000 218112 3052
rect 222660 3000 222712 3052
rect 225512 3000 225564 3052
rect 229284 3000 229336 3052
rect 229836 3000 229888 3052
rect 233700 3000 233752 3052
rect 234620 3000 234672 3052
rect 238116 3000 238168 3052
rect 240508 3000 240560 3052
rect 243636 3000 243688 3052
rect 248788 3000 248840 3052
rect 251364 3000 251416 3052
rect 331312 3000 331364 3052
rect 333888 3000 333940 3052
rect 334808 3000 334860 3052
rect 337476 3000 337528 3052
rect 513472 3000 513524 3052
rect 529020 3000 529072 3052
rect 535552 3000 535604 3052
rect 542820 3000 542872 3052
rect 543464 3000 543516 3052
rect 560484 3000 560536 3052
rect 564348 3000 564400 3052
rect 583392 3000 583444 3052
rect 203892 2932 203944 2984
rect 209412 2932 209464 2984
rect 212172 2932 212224 2984
rect 217140 2932 217192 2984
rect 222752 2932 222804 2984
rect 227352 2932 227404 2984
rect 227536 2932 227588 2984
rect 231768 2932 231820 2984
rect 232228 2932 232280 2984
rect 236184 2932 236236 2984
rect 237012 2932 237064 2984
rect 240600 2932 240652 2984
rect 242900 2932 242952 2984
rect 246120 2932 246172 2984
rect 246396 2932 246448 2984
rect 249432 2932 249484 2984
rect 253480 2932 253532 2984
rect 256056 2932 256108 2984
rect 310244 2932 310296 2984
rect 311440 2932 311492 2984
rect 325700 2932 325752 2984
rect 328000 2932 328052 2984
rect 329012 2932 329064 2984
rect 331588 2932 331640 2984
rect 332324 2932 332376 2984
rect 335084 2932 335136 2984
rect 341156 2932 341208 2984
rect 344560 2932 344612 2984
rect 514852 2932 514904 2984
rect 521844 2932 521896 2984
rect 536564 2932 536616 2984
rect 553768 2932 553820 2984
rect 148324 2864 148376 2916
rect 157524 2864 157576 2916
rect 157800 2864 157852 2916
rect 166632 2864 166684 2916
rect 169576 2864 169628 2916
rect 177672 2864 177724 2916
rect 177856 2864 177908 2916
rect 185400 2864 185452 2916
rect 99840 2796 99892 2848
rect 112260 2796 112312 2848
rect 118792 2796 118844 2848
rect 129648 2796 129700 2848
rect 132960 2796 133012 2848
rect 143448 2796 143500 2848
rect 150624 2796 150676 2848
rect 160008 2796 160060 2848
rect 161296 2796 161348 2848
rect 169944 2796 169996 2848
rect 170772 2796 170824 2848
rect 178776 2796 178828 2848
rect 180248 2796 180300 2848
rect 187608 2864 187660 2916
rect 192392 2864 192444 2916
rect 198372 2864 198424 2916
rect 199108 2864 199160 2916
rect 204996 2864 205048 2916
rect 205088 2864 205140 2916
rect 210516 2864 210568 2916
rect 213368 2864 213420 2916
rect 218244 2864 218296 2916
rect 219256 2864 219308 2916
rect 223488 2864 223540 2916
rect 223948 2864 224000 2916
rect 228456 2864 228508 2916
rect 228732 2864 228784 2916
rect 232872 2864 232924 2916
rect 235816 2864 235868 2916
rect 239496 2864 239548 2916
rect 242072 2864 242124 2916
rect 245016 2864 245068 2916
rect 245200 2864 245252 2916
rect 248328 2864 248380 2916
rect 249984 2864 250036 2916
rect 252744 2864 252796 2916
rect 254676 2864 254728 2916
rect 257160 2864 257212 2916
rect 261760 2864 261812 2916
rect 263784 2864 263836 2916
rect 312452 2864 312504 2916
rect 313832 2864 313884 2916
rect 314568 2864 314620 2916
rect 316224 2864 316276 2916
rect 316868 2864 316920 2916
rect 318524 2864 318576 2916
rect 319076 2864 319128 2916
rect 320916 2864 320968 2916
rect 321284 2864 321336 2916
rect 323308 2864 323360 2916
rect 323492 2864 323544 2916
rect 325608 2864 325660 2916
rect 327908 2864 327960 2916
rect 330392 2864 330444 2916
rect 333428 2864 333480 2916
rect 336280 2864 336332 2916
rect 340052 2864 340104 2916
rect 342996 2864 343048 2916
rect 514760 2864 514812 2916
rect 523040 2864 523092 2916
rect 525800 2864 525852 2916
rect 531320 2864 531372 2916
rect 532240 2864 532292 2916
rect 539600 2864 539652 2916
rect 187332 2796 187384 2848
rect 194232 2796 194284 2848
rect 194416 2796 194468 2848
rect 200856 2796 200908 2848
rect 202696 2796 202748 2848
rect 208400 2796 208452 2848
rect 208584 2796 208636 2848
rect 213828 2796 213880 2848
rect 215668 2796 215720 2848
rect 220728 2796 220780 2848
rect 221556 2796 221608 2848
rect 226248 2796 226300 2848
rect 226340 2796 226392 2848
rect 230664 2796 230716 2848
rect 233424 2796 233476 2848
rect 237288 2796 237340 2848
rect 238116 2796 238168 2848
rect 241704 2796 241756 2848
rect 244096 2796 244148 2848
rect 247224 2796 247276 2848
rect 247592 2796 247644 2848
rect 250536 2796 250588 2848
rect 252376 2796 252428 2848
rect 254952 2796 255004 2848
rect 255872 2796 255924 2848
rect 258264 2796 258316 2848
rect 260656 2796 260708 2848
rect 262680 2796 262732 2848
rect 304724 2796 304776 2848
rect 305552 2796 305604 2848
rect 306932 2796 306984 2848
rect 307944 2796 307996 2848
rect 309140 2796 309192 2848
rect 310244 2796 310296 2848
rect 311348 2796 311400 2848
rect 312636 2796 312688 2848
rect 313556 2796 313608 2848
rect 315028 2796 315080 2848
rect 315764 2796 315816 2848
rect 317328 2796 317380 2848
rect 317972 2796 318024 2848
rect 319720 2796 319772 2848
rect 320088 2796 320140 2848
rect 322112 2796 322164 2848
rect 322388 2796 322440 2848
rect 324412 2796 324464 2848
rect 324596 2796 324648 2848
rect 326804 2796 326856 2848
rect 326988 2796 327040 2848
rect 329196 2796 329248 2848
rect 330116 2796 330168 2848
rect 332692 2796 332744 2848
rect 335636 2796 335688 2848
rect 338672 2796 338724 2848
rect 338948 2796 339000 2848
rect 342076 2796 342128 2848
rect 346676 2796 346728 2848
rect 350448 2796 350500 2848
rect 353208 2796 353260 2848
rect 357532 2796 357584 2848
rect 372344 2796 372396 2848
rect 377680 2796 377732 2848
rect 520188 2796 520240 2848
rect 536840 2796 536892 2848
rect 541992 2864 542044 2916
rect 561956 2864 562008 2916
rect 581000 2864 581052 2916
rect 541532 2796 541584 2848
rect 550272 2796 550324 2848
rect 559748 2796 559800 2848
rect 578608 2796 578660 2848
rect 525432 2728 525484 2780
rect 77116 1300 77168 1352
rect 82728 1300 82780 1352
rect 88984 1300 89036 1352
rect 93768 1300 93820 1352
rect 95148 1300 95200 1352
rect 99288 1300 99340 1352
rect 198280 1300 198332 1352
rect 204168 1300 204220 1352
rect 207388 1300 207440 1352
rect 213000 1300 213052 1352
rect 257068 1300 257120 1352
rect 259368 1300 259420 1352
rect 259460 1300 259512 1352
rect 261576 1300 261628 1352
rect 262956 1300 263008 1352
rect 264888 1300 264940 1352
rect 265348 1300 265400 1352
rect 267096 1300 267148 1352
rect 267740 1300 267792 1352
rect 269304 1300 269356 1352
rect 271236 1300 271288 1352
rect 272616 1300 272668 1352
rect 273628 1300 273680 1352
rect 274824 1300 274876 1352
rect 277124 1300 277176 1352
rect 278136 1300 278188 1352
rect 279516 1300 279568 1352
rect 280344 1300 280396 1352
rect 336648 1300 336700 1352
rect 339868 1300 339920 1352
rect 342168 1300 342220 1352
rect 345756 1300 345808 1352
rect 348884 1300 348936 1352
rect 352840 1300 352892 1352
rect 356612 1300 356664 1352
rect 361120 1300 361172 1352
rect 364248 1300 364300 1352
rect 369400 1300 369452 1352
rect 374276 1300 374328 1352
rect 379612 1300 379664 1352
rect 385316 1300 385368 1352
rect 391848 1300 391900 1352
rect 396356 1300 396408 1352
rect 403624 1300 403676 1352
rect 406292 1300 406344 1352
rect 414296 1300 414348 1352
rect 415124 1300 415176 1352
rect 423404 1300 423456 1352
rect 428372 1300 428424 1352
rect 437572 1300 437624 1352
rect 439412 1300 439464 1352
rect 443736 1300 443788 1352
rect 85488 1232 85540 1284
rect 89352 1232 89404 1284
rect 92940 1232 92992 1284
rect 97080 1232 97132 1284
rect 258264 1232 258316 1284
rect 260472 1232 260524 1284
rect 264152 1232 264204 1284
rect 265992 1232 266044 1284
rect 266544 1232 266596 1284
rect 268200 1232 268252 1284
rect 270040 1232 270092 1284
rect 271512 1232 271564 1284
rect 272432 1232 272484 1284
rect 273720 1232 273772 1284
rect 343364 1232 343416 1284
rect 346952 1232 347004 1284
rect 349988 1232 350040 1284
rect 354036 1232 354088 1284
rect 357716 1232 357768 1284
rect 362316 1232 362368 1284
rect 365444 1232 365496 1284
rect 370228 1232 370280 1284
rect 370964 1232 371016 1284
rect 376116 1232 376168 1284
rect 376484 1232 376536 1284
rect 382372 1232 382424 1284
rect 388628 1232 388680 1284
rect 395344 1232 395396 1284
rect 404084 1232 404136 1284
rect 411904 1232 411956 1284
rect 413928 1232 413980 1284
rect 422576 1232 422628 1284
rect 426164 1232 426216 1284
rect 435180 1232 435232 1284
rect 436008 1232 436060 1284
rect 445852 1300 445904 1352
rect 449348 1300 449400 1352
rect 453212 1300 453264 1352
rect 444932 1232 444984 1284
rect 455696 1300 455748 1352
rect 462596 1300 462648 1352
rect 474188 1300 474240 1352
rect 475844 1300 475896 1352
rect 488816 1300 488868 1352
rect 493508 1300 493560 1352
rect 507308 1300 507360 1352
rect 526628 1300 526680 1352
rect 535552 1300 535604 1352
rect 539876 1300 539928 1352
rect 556988 1300 557040 1352
rect 454868 1232 454920 1284
rect 466000 1232 466052 1284
rect 469128 1232 469180 1284
rect 481364 1232 481416 1284
rect 495716 1232 495768 1284
rect 509700 1232 509752 1284
rect 510068 1232 510120 1284
rect 520188 1232 520240 1284
rect 524328 1232 524380 1284
rect 532608 1232 532660 1284
rect 68836 1164 68888 1216
rect 79416 1164 79468 1216
rect 268844 1164 268896 1216
rect 270408 1164 270460 1216
rect 359924 1164 359976 1216
rect 364616 1164 364668 1216
rect 368756 1164 368808 1216
rect 373908 1164 373960 1216
rect 378692 1164 378744 1216
rect 384396 1164 384448 1216
rect 387524 1164 387576 1216
rect 394240 1164 394292 1216
rect 395252 1164 395304 1216
rect 402520 1164 402572 1216
rect 420644 1164 420696 1216
rect 429292 1164 429344 1216
rect 434996 1164 435048 1216
rect 445024 1164 445076 1216
rect 352196 1096 352248 1148
rect 356336 1096 356388 1148
rect 361028 1096 361080 1148
rect 365444 1096 365496 1148
rect 369768 1096 369820 1148
rect 375288 1096 375340 1148
rect 379796 1096 379848 1148
rect 385960 1096 386012 1148
rect 397368 1096 397420 1148
rect 404820 1096 404872 1148
rect 412916 1096 412968 1148
rect 421380 1096 421432 1148
rect 422852 1096 422904 1148
rect 431868 1096 431920 1148
rect 438308 1096 438360 1148
rect 445760 1096 445812 1148
rect 355508 1028 355560 1080
rect 359924 1028 359976 1080
rect 366548 1028 366600 1080
rect 371332 1028 371384 1080
rect 373172 1028 373224 1080
rect 378508 1028 378560 1080
rect 394148 1028 394200 1080
rect 401324 1028 401376 1080
rect 424968 1028 425020 1080
rect 434076 1028 434128 1080
rect 442724 1028 442776 1080
rect 450452 1164 450504 1216
rect 461584 1164 461636 1216
rect 482468 1164 482520 1216
rect 495532 1164 495584 1216
rect 506756 1164 506808 1216
rect 514852 1164 514904 1216
rect 528836 1164 528888 1216
rect 545488 1164 545540 1216
rect 453304 1096 453356 1148
rect 455972 1096 456024 1148
rect 467472 1096 467524 1148
rect 474648 1096 474700 1148
rect 487252 1096 487304 1148
rect 487988 1096 488040 1148
rect 501420 1096 501472 1148
rect 507768 1096 507820 1148
rect 514760 1096 514812 1148
rect 533252 1096 533304 1148
rect 541532 1096 541584 1148
rect 446036 1028 446088 1080
rect 345572 960 345624 1012
rect 349252 960 349304 1012
rect 351092 960 351144 1012
rect 355232 960 355284 1012
rect 362132 960 362184 1012
rect 367008 960 367060 1012
rect 367652 960 367704 1012
rect 372896 960 372948 1012
rect 375196 960 375248 1012
rect 381176 960 381228 1012
rect 419448 960 419500 1012
rect 428464 960 428516 1012
rect 431684 960 431736 1012
rect 441436 960 441488 1012
rect 441528 960 441580 1012
rect 448520 960 448572 1012
rect 19432 892 19484 944
rect 37464 892 37516 944
rect 358728 892 358780 944
rect 363512 892 363564 944
rect 377588 892 377640 944
rect 383568 892 383620 944
rect 416228 892 416280 944
rect 424968 892 425020 944
rect 430488 892 430540 944
rect 21824 824 21876 876
rect 39672 824 39724 876
rect 337844 824 337896 876
rect 340972 824 341024 876
rect 347688 824 347740 876
rect 351644 824 351696 876
rect 386328 824 386380 876
rect 392676 824 392728 876
rect 421748 824 421800 876
rect 430856 824 430908 876
rect 437204 892 437256 944
rect 447416 892 447468 944
rect 451556 1028 451608 1080
rect 462412 1028 462464 1080
rect 485688 1028 485740 1080
rect 490104 1028 490156 1080
rect 490196 1028 490248 1080
rect 494796 1028 494848 1080
rect 525524 1028 525576 1080
rect 536840 1028 536892 1080
rect 448704 960 448756 1012
rect 451740 960 451792 1012
rect 453212 960 453264 1012
rect 456892 892 456944 944
rect 457076 960 457128 1012
rect 468300 960 468352 1012
rect 486884 960 486936 1012
rect 500592 960 500644 1012
rect 501236 960 501288 1012
rect 515496 960 515548 1012
rect 515588 960 515640 1012
rect 525800 960 525852 1012
rect 527732 960 527784 1012
rect 544384 960 544436 1012
rect 460020 892 460072 944
rect 481548 892 481600 944
rect 440332 824 440384 876
rect 447048 824 447100 876
rect 458088 824 458140 876
rect 494612 892 494664 944
rect 508872 892 508924 944
rect 520004 892 520056 944
rect 536104 892 536156 944
rect 494704 824 494756 876
rect 494796 824 494848 876
rect 503812 824 503864 876
rect 523316 824 523368 876
rect 532240 824 532292 876
rect 547604 824 547656 876
rect 565636 824 565688 876
rect 8760 756 8812 808
rect 27528 756 27580 808
rect 251180 756 251232 808
rect 253848 756 253900 808
rect 429476 756 429528 808
rect 439136 756 439188 808
rect 440516 756 440568 808
rect 450912 756 450964 808
rect 483572 756 483624 808
rect 497096 756 497148 808
rect 514484 756 514536 808
rect 529756 756 529808 808
rect 532148 756 532200 808
rect 548708 756 548760 808
rect 550916 756 550968 808
rect 569132 756 569184 808
rect 17040 688 17092 740
rect 35256 688 35308 740
rect 432788 688 432840 740
rect 442632 688 442684 740
rect 443828 688 443880 740
rect 454132 688 454184 740
rect 468116 688 468168 740
rect 480536 688 480588 740
rect 489092 688 489144 740
rect 502984 688 503036 740
rect 522212 688 522264 740
rect 538220 688 538272 740
rect 540888 688 540940 740
rect 558552 688 558604 740
rect 15936 620 15988 672
rect 34152 620 34204 672
rect 35992 620 36044 672
rect 52920 620 52972 672
rect 11152 552 11204 604
rect 29736 552 29788 604
rect 39580 552 39632 604
rect 56232 552 56284 604
rect 384212 552 384264 604
rect 390652 552 390704 604
rect 393044 552 393096 604
rect 400128 620 400180 672
rect 401876 620 401928 672
rect 409236 620 409288 672
rect 397736 552 397788 604
rect 408408 552 408460 604
rect 409604 552 409656 604
rect 417884 620 417936 672
rect 427268 620 427320 672
rect 436744 620 436796 672
rect 448244 620 448296 672
rect 459192 620 459244 672
rect 459284 620 459336 672
rect 471060 620 471112 672
rect 471428 620 471480 672
rect 479524 620 479576 672
rect 480168 620 480220 672
rect 493140 620 493192 672
rect 502248 620 502300 672
rect 517152 620 517204 672
rect 542084 620 542136 672
rect 559748 620 559800 672
rect 416688 552 416740 604
rect 433892 552 433944 604
rect 443460 552 443512 604
rect 443736 552 443788 604
rect 449808 552 449860 604
rect 461492 552 461544 604
rect 473452 552 473504 604
rect 491208 552 491260 604
rect 505376 552 505428 604
rect 508964 552 509016 604
rect 524236 552 524288 604
rect 545396 552 545448 604
rect 563244 620 563296 672
rect 562048 552 562100 604
rect 18052 484 18104 536
rect 36360 484 36412 536
rect 38568 484 38620 536
rect 55128 484 55180 536
rect 390836 484 390888 536
rect 14556 416 14608 468
rect 33048 416 33100 468
rect 34612 416 34664 468
rect 51816 416 51868 468
rect 382004 416 382056 468
rect 387892 416 387944 468
rect 470324 484 470376 536
rect 482468 484 482520 536
rect 490104 484 490156 536
rect 499120 484 499172 536
rect 503444 484 503496 536
rect 517980 484 518032 536
rect 544568 484 544620 536
rect 464804 416 464856 468
rect 476580 416 476632 468
rect 478328 416 478380 468
rect 490748 416 490800 468
rect 497924 416 497976 468
rect 512092 416 512144 468
rect 516692 416 516744 468
rect 532148 416 532200 468
rect 548892 416 548944 468
rect 567016 416 567068 468
rect 9772 348 9824 400
rect 28632 348 28684 400
rect 32220 348 32272 400
rect 49608 348 49660 400
rect 405188 348 405240 400
rect 412824 348 412876 400
rect 418436 348 418488 400
rect 426900 348 426952 400
rect 453764 348 453816 400
rect 464988 348 465040 400
rect 472532 348 472584 400
rect 3240 280 3292 332
rect 22008 280 22060 332
rect 22836 280 22888 332
rect 40500 280 40552 332
rect 42892 280 42944 332
rect 59360 280 59412 332
rect 391664 280 391716 332
rect 398748 280 398800 332
rect 400772 280 400824 332
rect 408592 280 408644 332
rect 412088 280 412140 332
rect 420368 280 420420 332
rect 457904 280 457956 332
rect 470048 280 470100 332
rect 479156 280 479208 332
rect 479524 348 479576 400
rect 484216 348 484268 400
rect 499028 348 499080 400
rect 513380 348 513432 400
rect 517796 348 517848 400
rect 533896 348 533948 400
rect 534356 348 534408 400
rect 551100 348 551152 400
rect 555332 348 555384 400
rect 573548 348 573600 400
rect 484860 280 484912 332
rect 504548 280 504600 332
rect 519728 280 519780 332
rect 521108 280 521160 332
rect 537392 280 537444 332
rect 538772 280 538824 332
rect 556344 280 556396 332
rect 557172 280 557224 332
rect 575940 280 575992 332
rect 3884 212 3936 264
rect 23204 212 23256 264
rect 24584 212 24636 264
rect 41604 212 41656 264
rect 42248 212 42300 264
rect 58164 212 58216 264
rect 380808 212 380860 264
rect 386788 212 386840 264
rect 398564 212 398616 264
rect 406200 212 406252 264
rect 410984 212 411036 264
rect 418620 212 418672 264
rect 445760 212 445812 264
rect 448244 212 448296 264
rect 465908 212 465960 264
rect 478328 212 478380 264
rect 492496 212 492548 264
rect 492588 212 492640 264
rect 506664 212 506716 264
rect 511448 212 511500 264
rect 526260 212 526312 264
rect 535368 212 535420 264
rect 552848 212 552900 264
rect 554228 212 554280 264
rect 572904 212 572956 264
rect 8024 144 8076 196
rect 26332 144 26384 196
rect 30288 144 30340 196
rect 47400 144 47452 196
rect 389732 144 389784 196
rect 396172 144 396224 196
rect 399668 144 399720 196
rect 407028 144 407080 196
rect 407396 144 407448 196
rect 415308 144 415360 196
rect 417332 144 417384 196
rect 425796 144 425848 196
rect 452568 144 452620 196
rect 464160 144 464212 196
rect 467012 144 467064 196
rect 478972 144 479024 196
rect 484676 144 484728 196
rect 498384 144 498436 196
rect 505652 144 505704 196
rect 520372 144 520424 196
rect 537668 144 537720 196
rect 554780 144 554832 196
rect 558828 144 558880 196
rect 577136 144 577188 196
rect 1492 76 1544 128
rect 20904 76 20956 128
rect 31116 76 31168 128
rect 48504 76 48556 128
rect 53564 76 53616 128
rect 69480 76 69532 128
rect 354404 76 354456 128
rect 358912 76 358964 128
rect 363236 76 363288 128
rect 367836 76 367888 128
rect 402888 76 402940 128
rect 410984 76 411036 128
rect 460664 76 460716 128
rect 472440 76 472492 128
rect 473636 76 473688 128
rect 486608 76 486660 128
rect 500132 76 500184 128
rect 514944 76 514996 128
rect 518808 76 518860 128
rect 534540 76 534592 128
rect 546408 76 546460 128
rect 564624 76 564676 128
rect 388 8 440 60
rect 19800 8 19852 60
rect 20444 8 20496 60
rect 38200 8 38252 60
rect 45284 8 45336 60
rect 61752 8 61804 60
rect 344744 8 344796 60
rect 348240 8 348292 60
rect 383108 8 383160 60
rect 389640 8 389692 60
rect 423956 8 424008 60
rect 433432 8 433484 60
rect 463608 8 463660 60
rect 475936 8 475988 60
rect 477224 8 477276 60
rect 490104 8 490156 60
rect 496728 8 496780 60
rect 511448 8 511500 60
rect 512644 8 512696 60
rect 528008 8 528060 60
rect 531044 8 531096 60
rect 548064 8 548116 60
rect 551928 8 551980 60
rect 570512 8 570564 60
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 251652 703582 251864 703610
rect 8128 701010 8156 703520
rect 24320 702506 24348 703520
rect 24308 702500 24360 702506
rect 24308 702442 24360 702448
rect 29276 702500 29328 702506
rect 29276 702442 29328 702448
rect 8116 701004 8168 701010
rect 8116 700946 8168 700952
rect 13084 701004 13136 701010
rect 13084 700946 13136 700952
rect 13096 700890 13124 700946
rect 13096 700862 13386 700890
rect 29288 700876 29316 702442
rect 40512 701010 40540 703520
rect 56796 701010 56824 703520
rect 72988 701010 73016 703520
rect 89180 701010 89208 703520
rect 105464 701010 105492 703520
rect 121656 701010 121684 703520
rect 137848 701010 137876 703520
rect 154132 701010 154160 703520
rect 170324 701010 170352 703520
rect 186516 703050 186544 703520
rect 186504 703044 186556 703050
rect 186504 702986 186556 702992
rect 188436 703044 188488 703050
rect 188436 702986 188488 702992
rect 40500 701004 40552 701010
rect 40500 700946 40552 700952
rect 44916 701004 44968 701010
rect 44916 700946 44968 700952
rect 56784 701004 56836 701010
rect 56784 700946 56836 700952
rect 60740 701004 60792 701010
rect 60740 700946 60792 700952
rect 72976 701004 73028 701010
rect 72976 700946 73028 700952
rect 76748 701004 76800 701010
rect 76748 700946 76800 700952
rect 89168 701004 89220 701010
rect 89168 700946 89220 700952
rect 92572 701004 92624 701010
rect 92572 700946 92624 700952
rect 105452 701004 105504 701010
rect 105452 700946 105504 700952
rect 108580 701004 108632 701010
rect 108580 700946 108632 700952
rect 121644 701004 121696 701010
rect 121644 700946 121696 700952
rect 124404 701004 124456 701010
rect 124404 700946 124456 700952
rect 137836 701004 137888 701010
rect 137836 700946 137888 700952
rect 140412 701004 140464 701010
rect 140412 700946 140464 700952
rect 154120 701004 154172 701010
rect 154120 700946 154172 700952
rect 156236 701004 156288 701010
rect 156236 700946 156288 700952
rect 170312 701004 170364 701010
rect 170312 700946 170364 700952
rect 172428 701004 172480 701010
rect 172428 700946 172480 700952
rect 44928 700890 44956 700946
rect 60752 700890 60780 700946
rect 76760 700890 76788 700946
rect 92584 700890 92612 700946
rect 108592 700890 108620 700946
rect 124416 700890 124444 700946
rect 140424 700890 140452 700946
rect 156248 700890 156276 700946
rect 172440 700890 172468 700946
rect 44928 700862 45218 700890
rect 60752 700862 61134 700890
rect 76760 700862 77050 700890
rect 92584 700862 92966 700890
rect 108592 700862 108882 700890
rect 124416 700862 124798 700890
rect 140424 700862 140714 700890
rect 156248 700862 156630 700890
rect 172440 700862 172546 700890
rect 188448 700876 188476 702986
rect 202800 701010 202828 703520
rect 218992 702506 219020 703520
rect 235184 703050 235212 703520
rect 251468 703474 251496 703520
rect 251652 703474 251680 703582
rect 251468 703446 251680 703474
rect 235172 703044 235224 703050
rect 235172 702986 235224 702992
rect 236184 703044 236236 703050
rect 236184 702986 236236 702992
rect 218980 702500 219032 702506
rect 218980 702442 219032 702448
rect 220268 702500 220320 702506
rect 220268 702442 220320 702448
rect 202788 701004 202840 701010
rect 202788 700946 202840 700952
rect 204260 701004 204312 701010
rect 204260 700946 204312 700952
rect 204272 700890 204300 700946
rect 204272 700862 204378 700890
rect 220280 700876 220308 702442
rect 236196 700876 236224 702986
rect 251836 700890 251864 703582
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332152 703582 332364 703610
rect 267660 700890 267688 703520
rect 283852 700890 283880 703520
rect 300136 700890 300164 703520
rect 316328 702434 316356 703520
rect 316052 702406 316356 702434
rect 316052 700890 316080 702406
rect 332152 700890 332180 703582
rect 332336 703474 332364 703582
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 332520 703474 332548 703520
rect 332336 703446 332548 703474
rect 348804 701010 348832 703520
rect 364996 701010 365024 703520
rect 381188 701010 381216 703520
rect 397472 701010 397500 703520
rect 413664 701010 413692 703520
rect 429856 701010 429884 703520
rect 446140 701010 446168 703520
rect 462332 702506 462360 703520
rect 459100 702500 459152 702506
rect 459100 702442 459152 702448
rect 462320 702500 462372 702506
rect 462320 702442 462372 702448
rect 348056 701004 348108 701010
rect 348056 700946 348108 700952
rect 348792 701004 348844 701010
rect 348792 700946 348844 700952
rect 363880 701004 363932 701010
rect 363880 700946 363932 700952
rect 364984 701004 365036 701010
rect 364984 700946 365036 700952
rect 379336 701004 379388 701010
rect 379336 700946 379388 700952
rect 381176 701004 381228 701010
rect 381176 700946 381228 700952
rect 395712 701004 395764 701010
rect 395712 700946 395764 700952
rect 397460 701004 397512 701010
rect 397460 700946 397512 700952
rect 411720 701004 411772 701010
rect 411720 700946 411772 700952
rect 413652 701004 413704 701010
rect 413652 700946 413704 700952
rect 427544 701004 427596 701010
rect 427544 700946 427596 700952
rect 429844 701004 429896 701010
rect 429844 700946 429896 700952
rect 443552 701004 443604 701010
rect 443552 700946 443604 700952
rect 446128 701004 446180 701010
rect 446128 700946 446180 700952
rect 348068 700890 348096 700946
rect 363892 700890 363920 700946
rect 251836 700862 252126 700890
rect 267660 700862 268042 700890
rect 283852 700862 283958 700890
rect 299966 700862 300164 700890
rect 315882 700862 316080 700890
rect 331798 700862 332180 700890
rect 347714 700862 348096 700890
rect 363630 700862 363920 700890
rect 379348 700890 379376 700946
rect 395724 700890 395752 700946
rect 411732 700890 411760 700946
rect 427556 700890 427584 700946
rect 443564 700890 443592 700946
rect 379348 700862 379454 700890
rect 395462 700862 395752 700890
rect 411378 700862 411760 700890
rect 427294 700862 427584 700890
rect 443210 700862 443592 700890
rect 459112 700876 459140 702442
rect 478524 701010 478552 703520
rect 494808 702778 494836 703520
rect 490932 702772 490984 702778
rect 490932 702714 490984 702720
rect 494796 702772 494848 702778
rect 494796 702714 494848 702720
rect 475384 701004 475436 701010
rect 475384 700946 475436 700952
rect 478512 701004 478564 701010
rect 478512 700946 478564 700952
rect 475396 700890 475424 700946
rect 475042 700862 475424 700890
rect 490944 700876 490972 702714
rect 511000 702506 511028 703520
rect 527192 703066 527220 703520
rect 527100 703050 527220 703066
rect 522764 703044 522816 703050
rect 522764 702986 522816 702992
rect 527088 703044 527220 703050
rect 527140 703038 527220 703044
rect 527088 702986 527140 702992
rect 506848 702500 506900 702506
rect 506848 702442 506900 702448
rect 510988 702500 511040 702506
rect 510988 702442 511040 702448
rect 506860 700876 506888 702442
rect 522776 700876 522804 702986
rect 543476 702778 543504 703520
rect 538680 702772 538732 702778
rect 538680 702714 538732 702720
rect 543464 702772 543516 702778
rect 543464 702714 543516 702720
rect 538692 700876 538720 702714
rect 559668 702506 559696 703520
rect 575860 703050 575888 703520
rect 570512 703044 570564 703050
rect 570512 702986 570564 702992
rect 575848 703044 575900 703050
rect 575848 702986 575900 702992
rect 554596 702500 554648 702506
rect 554596 702442 554648 702448
rect 559656 702500 559708 702506
rect 559656 702442 559708 702448
rect 554608 700876 554636 702442
rect 570524 700876 570552 702986
rect 2778 697368 2834 697377
rect 2778 697303 2834 697312
rect 2792 690849 2820 697303
rect 581642 697232 581698 697241
rect 581642 697167 581698 697176
rect 581656 691529 581684 697167
rect 581642 691520 581698 691529
rect 581642 691455 581698 691464
rect 2778 690840 2834 690849
rect 2778 690775 2834 690784
rect 2778 684312 2834 684321
rect 2778 684247 2834 684256
rect 2792 678065 2820 684247
rect 582378 683904 582434 683913
rect 582378 683839 582434 683848
rect 582392 678473 582420 683839
rect 582378 678464 582434 678473
rect 582378 678399 582434 678408
rect 2778 678056 2834 678065
rect 2778 677991 2834 678000
rect 2778 671256 2834 671265
rect 2778 671191 2834 671200
rect 2792 665281 2820 671191
rect 582378 670712 582434 670721
rect 582378 670647 582434 670656
rect 582392 665417 582420 670647
rect 582378 665408 582434 665417
rect 582378 665343 582434 665352
rect 2778 665272 2834 665281
rect 2778 665207 2834 665216
rect 2778 658200 2834 658209
rect 2778 658135 2834 658144
rect 2792 652497 2820 658135
rect 582378 657384 582434 657393
rect 582378 657319 582434 657328
rect 2778 652488 2834 652497
rect 2778 652423 2834 652432
rect 582392 652361 582420 657319
rect 582378 652352 582434 652361
rect 582378 652287 582434 652296
rect 2778 645144 2834 645153
rect 2778 645079 2834 645088
rect 2792 639713 2820 645079
rect 581642 644056 581698 644065
rect 581642 643991 581698 644000
rect 2778 639704 2834 639713
rect 2778 639639 2834 639648
rect 581656 639305 581684 643991
rect 581642 639296 581698 639305
rect 581642 639231 581698 639240
rect 2778 632088 2834 632097
rect 2778 632023 2834 632032
rect 2792 626929 2820 632023
rect 582378 630864 582434 630873
rect 582378 630799 582434 630808
rect 2778 626920 2834 626929
rect 2778 626855 2834 626864
rect 582392 626249 582420 630799
rect 582378 626240 582434 626249
rect 582378 626175 582434 626184
rect 2778 619168 2834 619177
rect 2778 619103 2834 619112
rect 2792 614009 2820 619103
rect 581642 617536 581698 617545
rect 581642 617471 581698 617480
rect 2778 614000 2834 614009
rect 2778 613935 2834 613944
rect 581656 613193 581684 617471
rect 581642 613184 581698 613193
rect 581642 613119 581698 613128
rect 2778 606112 2834 606121
rect 2778 606047 2834 606056
rect 2792 601361 2820 606047
rect 581642 604208 581698 604217
rect 581642 604143 581698 604152
rect 2778 601352 2834 601361
rect 2778 601287 2834 601296
rect 581656 600137 581684 604143
rect 581642 600128 581698 600137
rect 581642 600063 581698 600072
rect 1582 593056 1638 593065
rect 1582 592991 1638 593000
rect 1596 588577 1624 592991
rect 581642 591016 581698 591025
rect 581642 590951 581698 590960
rect 1582 588568 1638 588577
rect 1582 588503 1638 588512
rect 581656 587081 581684 590951
rect 581642 587072 581698 587081
rect 581642 587007 581698 587016
rect 2042 580000 2098 580009
rect 2042 579935 2098 579944
rect 2056 575793 2084 579935
rect 581642 577688 581698 577697
rect 581642 577623 581698 577632
rect 2042 575784 2098 575793
rect 2042 575719 2098 575728
rect 581656 574025 581684 577623
rect 581642 574016 581698 574025
rect 581642 573951 581698 573960
rect 1490 566944 1546 566953
rect 1490 566879 1546 566888
rect 1504 563009 1532 566879
rect 582378 564360 582434 564369
rect 582378 564295 582434 564304
rect 1490 563000 1546 563009
rect 1490 562935 1546 562944
rect 582392 560969 582420 564295
rect 582378 560960 582434 560969
rect 582378 560895 582434 560904
rect 1490 553888 1546 553897
rect 1490 553823 1546 553832
rect 1504 550225 1532 553823
rect 581642 551168 581698 551177
rect 581642 551103 581698 551112
rect 1490 550216 1546 550225
rect 1490 550151 1546 550160
rect 581656 547777 581684 551103
rect 581642 547768 581698 547777
rect 581642 547703 581698 547712
rect 1398 540832 1454 540841
rect 1398 540767 1454 540776
rect 1412 537441 1440 540767
rect 582378 537840 582434 537849
rect 582378 537775 582434 537784
rect 1398 537432 1454 537441
rect 1398 537367 1454 537376
rect 582392 534857 582420 537775
rect 582378 534848 582434 534857
rect 582378 534783 582434 534792
rect 1490 527912 1546 527921
rect 1490 527847 1546 527856
rect 1504 524657 1532 527847
rect 1490 524648 1546 524657
rect 1490 524583 1546 524592
rect 582378 524512 582434 524521
rect 582378 524447 582434 524456
rect 582392 521801 582420 524447
rect 582378 521792 582434 521801
rect 582378 521727 582434 521736
rect 1582 514856 1638 514865
rect 1582 514791 1638 514800
rect 1596 511873 1624 514791
rect 1582 511864 1638 511873
rect 1582 511799 1638 511808
rect 582378 511320 582434 511329
rect 582378 511255 582434 511264
rect 582392 508745 582420 511255
rect 582378 508736 582434 508745
rect 582378 508671 582434 508680
rect 1582 501800 1638 501809
rect 1582 501735 1638 501744
rect 1596 499089 1624 501735
rect 1582 499080 1638 499089
rect 1582 499015 1638 499024
rect 581642 497992 581698 498001
rect 581642 497927 581698 497936
rect 581656 495689 581684 497927
rect 581642 495680 581698 495689
rect 581642 495615 581698 495624
rect 1582 488744 1638 488753
rect 1582 488679 1638 488688
rect 1596 486305 1624 488679
rect 1582 486296 1638 486305
rect 1582 486231 1638 486240
rect 582378 484664 582434 484673
rect 582378 484599 582434 484608
rect 582392 482633 582420 484599
rect 582378 482624 582434 482633
rect 582378 482559 582434 482568
rect 2778 475688 2834 475697
rect 2778 475623 2834 475632
rect 2792 473521 2820 475623
rect 2778 473512 2834 473521
rect 2778 473447 2834 473456
rect 581642 471472 581698 471481
rect 581642 471407 581698 471416
rect 581656 469577 581684 471407
rect 581642 469568 581698 469577
rect 581642 469503 581698 469512
rect 1582 462632 1638 462641
rect 1582 462567 1638 462576
rect 1596 460737 1624 462567
rect 1582 460728 1638 460737
rect 1582 460663 1638 460672
rect 581642 458144 581698 458153
rect 581642 458079 581698 458088
rect 581656 456521 581684 458079
rect 581642 456512 581698 456521
rect 581642 456447 581698 456456
rect 2778 449576 2834 449585
rect 2778 449511 2834 449520
rect 2792 447953 2820 449511
rect 2778 447944 2834 447953
rect 2778 447879 2834 447888
rect 2778 436656 2834 436665
rect 2778 436591 2834 436600
rect 2792 435169 2820 436591
rect 2778 435160 2834 435169
rect 2778 435095 2834 435104
rect 2778 423600 2834 423609
rect 2778 423535 2834 423544
rect 2792 422385 2820 423535
rect 2778 422376 2834 422385
rect 2778 422311 2834 422320
rect 1306 294400 1362 294409
rect 1306 294335 1362 294344
rect 1320 293185 1348 294335
rect 1306 293176 1362 293185
rect 1306 293111 1362 293120
rect 2778 281616 2834 281625
rect 2778 281551 2834 281560
rect 2792 280129 2820 281551
rect 2778 280120 2834 280129
rect 2778 280055 2834 280064
rect 1306 268832 1362 268841
rect 1306 268767 1362 268776
rect 1320 267209 1348 268767
rect 1306 267200 1362 267209
rect 1306 267135 1362 267144
rect 582378 260536 582434 260545
rect 582378 260471 582434 260480
rect 582392 258913 582420 260471
rect 582378 258904 582434 258913
rect 582378 258839 582434 258848
rect 1306 256048 1362 256057
rect 1306 255983 1362 255992
rect 1320 254153 1348 255983
rect 1306 254144 1362 254153
rect 1306 254079 1362 254088
rect 580906 247072 580962 247081
rect 580906 247007 580962 247016
rect 580920 245585 580948 247007
rect 580906 245576 580962 245585
rect 580906 245511 580962 245520
rect 2778 243264 2834 243273
rect 2778 243199 2834 243208
rect 2792 241097 2820 243199
rect 2778 241088 2834 241097
rect 2778 241023 2834 241032
rect 582378 234424 582434 234433
rect 582378 234359 582434 234368
rect 582392 232393 582420 234359
rect 582378 232384 582434 232393
rect 582378 232319 582434 232328
rect 2778 230616 2834 230625
rect 2778 230551 2834 230560
rect 2792 228041 2820 230551
rect 2778 228032 2834 228041
rect 2778 227967 2834 227976
rect 580906 220960 580962 220969
rect 580906 220895 580962 220904
rect 580920 219065 580948 220895
rect 580906 219056 580962 219065
rect 580906 218991 580962 219000
rect 2778 217696 2834 217705
rect 2778 217631 2834 217640
rect 2792 214985 2820 217631
rect 2778 214976 2834 214985
rect 2778 214911 2834 214920
rect 582378 208312 582434 208321
rect 582378 208247 582434 208256
rect 582392 205737 582420 208247
rect 582378 205728 582434 205737
rect 582378 205663 582434 205672
rect 2778 204912 2834 204921
rect 2778 204847 2834 204856
rect 2792 201929 2820 204847
rect 2778 201920 2834 201929
rect 2778 201855 2834 201864
rect 580906 194712 580962 194721
rect 580906 194647 580962 194656
rect 580920 192545 580948 194647
rect 580906 192536 580962 192545
rect 580906 192471 580962 192480
rect 1306 192128 1362 192137
rect 1306 192063 1362 192072
rect 1320 188873 1348 192063
rect 1306 188864 1362 188873
rect 1306 188799 1362 188808
rect 580906 182472 580962 182481
rect 580906 182407 580962 182416
rect 2778 179344 2834 179353
rect 2778 179279 2834 179288
rect 2792 175953 2820 179279
rect 580920 179217 580948 182407
rect 580906 179208 580962 179217
rect 580906 179143 580962 179152
rect 2778 175944 2834 175953
rect 2778 175879 2834 175888
rect 580906 168600 580962 168609
rect 580906 168535 580962 168544
rect 2778 166560 2834 166569
rect 2778 166495 2834 166504
rect 2792 162897 2820 166495
rect 580920 165889 580948 168535
rect 580906 165880 580962 165889
rect 580906 165815 580962 165824
rect 2778 162888 2834 162897
rect 2778 162823 2834 162832
rect 580906 156360 580962 156369
rect 580906 156295 580962 156304
rect 1306 153776 1362 153785
rect 1306 153711 1362 153720
rect 1320 149841 1348 153711
rect 580920 152697 580948 156295
rect 580906 152688 580962 152697
rect 580906 152623 580962 152632
rect 1306 149832 1362 149841
rect 1306 149767 1362 149776
rect 580906 142624 580962 142633
rect 580906 142559 580962 142568
rect 570 140992 626 141001
rect 570 140927 626 140936
rect 584 136785 612 140927
rect 580920 139369 580948 142559
rect 580906 139360 580962 139369
rect 580906 139295 580962 139304
rect 570 136776 626 136785
rect 570 136711 626 136720
rect 580906 130248 580962 130257
rect 580906 130183 580962 130192
rect 754 128208 810 128217
rect 754 128143 810 128152
rect 768 123729 796 128143
rect 580920 126041 580948 130183
rect 580906 126032 580962 126041
rect 580906 125967 580962 125976
rect 754 123720 810 123729
rect 754 123655 810 123664
rect 579894 116376 579950 116385
rect 579894 116311 579950 116320
rect 1306 115424 1362 115433
rect 1306 115359 1362 115368
rect 1320 110673 1348 115359
rect 579908 112849 579936 116311
rect 579894 112840 579950 112849
rect 579894 112775 579950 112784
rect 1306 110664 1362 110673
rect 1306 110599 1362 110608
rect 580906 103592 580962 103601
rect 580906 103527 580962 103536
rect 1582 102640 1638 102649
rect 1582 102575 1638 102584
rect 1596 97617 1624 102575
rect 580920 99521 580948 103527
rect 580906 99512 580962 99521
rect 580906 99447 580962 99456
rect 1582 97608 1638 97617
rect 1582 97543 1638 97552
rect 580906 90264 580962 90273
rect 580906 90199 580962 90208
rect 1582 89856 1638 89865
rect 1582 89791 1638 89800
rect 1596 84697 1624 89791
rect 580920 86193 580948 90199
rect 580906 86184 580962 86193
rect 580906 86119 580962 86128
rect 1582 84688 1638 84697
rect 1582 84623 1638 84632
rect 579894 77344 579950 77353
rect 579894 77279 579950 77288
rect 1582 77072 1638 77081
rect 1582 77007 1638 77016
rect 1596 71641 1624 77007
rect 579908 73001 579936 77279
rect 579894 72992 579950 73001
rect 579894 72927 579950 72936
rect 1582 71632 1638 71641
rect 1582 71567 1638 71576
rect 1490 64288 1546 64297
rect 1490 64223 1546 64232
rect 1504 58585 1532 64223
rect 580906 64152 580962 64161
rect 580906 64087 580962 64096
rect 580920 59673 580948 64087
rect 580906 59664 580962 59673
rect 580906 59599 580962 59608
rect 1490 58576 1546 58585
rect 1490 58511 1546 58520
rect 2042 51504 2098 51513
rect 2042 51439 2098 51448
rect 2056 45529 2084 51439
rect 580906 51096 580962 51105
rect 580906 51031 580962 51040
rect 580920 46345 580948 51031
rect 580906 46336 580962 46345
rect 580906 46271 580962 46280
rect 2042 45520 2098 45529
rect 2042 45455 2098 45464
rect 2042 38720 2098 38729
rect 2042 38655 2098 38664
rect 2056 32473 2084 38655
rect 580906 38040 580962 38049
rect 580906 37975 580962 37984
rect 580920 33153 580948 37975
rect 580906 33144 580962 33153
rect 580906 33079 580962 33088
rect 2042 32464 2098 32473
rect 2042 32399 2098 32408
rect 1490 25936 1546 25945
rect 1490 25871 1546 25880
rect 1504 19417 1532 25871
rect 580906 24984 580962 24993
rect 580906 24919 580962 24928
rect 580920 19825 580948 24919
rect 580906 19816 580962 19825
rect 580906 19751 580962 19760
rect 1490 19408 1546 19417
rect 1490 19343 1546 19352
rect 2042 13152 2098 13161
rect 2042 13087 2098 13096
rect 2056 6497 2084 13087
rect 582378 12472 582434 12481
rect 582378 12407 582434 12416
rect 582392 6633 582420 12407
rect 582378 6624 582434 6633
rect 582378 6559 582434 6568
rect 2042 6488 2098 6497
rect 2042 6423 2098 6432
rect 80256 3874 80546 3890
rect 101232 3874 101522 3890
rect 65524 3868 65576 3874
rect 65524 3810 65576 3816
rect 80244 3868 80546 3874
rect 80296 3862 80546 3868
rect 97632 3868 97684 3874
rect 80244 3810 80296 3816
rect 97632 3810 97684 3816
rect 101220 3868 101522 3874
rect 101272 3862 101522 3868
rect 101220 3810 101272 3816
rect 56048 3800 56100 3806
rect 56048 3742 56100 3748
rect 52552 3732 52604 3738
rect 52552 3674 52604 3680
rect 48964 3664 49016 3670
rect 48964 3606 49016 3612
rect 40960 3120 41012 3126
rect 19432 944 19484 950
rect 19432 886 19484 892
rect 8760 808 8812 814
rect 8760 750 8812 756
rect 8772 480 8800 750
rect 17040 740 17092 746
rect 17040 682 17092 688
rect 15936 672 15988 678
rect 15936 614 15988 620
rect 11152 604 11204 610
rect 11152 546 11204 552
rect 11164 480 11192 546
rect 12162 504 12218 513
rect 542 82 654 480
rect 400 66 654 82
rect 1492 128 1544 134
rect 1646 82 1758 480
rect 1544 76 1758 82
rect 1492 70 1758 76
rect 388 60 654 66
rect 440 54 654 60
rect 1504 54 1758 70
rect 388 2 440 8
rect 542 -960 654 54
rect 1646 -960 1758 54
rect 2842 354 2954 480
rect 2842 338 3280 354
rect 2842 332 3292 338
rect 2842 326 3240 332
rect 2842 -960 2954 326
rect 3240 274 3292 280
rect 3884 264 3936 270
rect 4038 218 4150 480
rect 3936 212 4150 218
rect 3884 206 4150 212
rect 3896 190 4150 206
rect 4038 -960 4150 190
rect 5234 82 5346 480
rect 6274 232 6330 241
rect 6430 218 6542 480
rect 6330 190 6542 218
rect 6274 167 6330 176
rect 5446 96 5502 105
rect 5234 54 5446 82
rect 5234 -960 5346 54
rect 5446 31 5502 40
rect 6430 -960 6542 190
rect 7626 218 7738 480
rect 7626 202 8064 218
rect 7626 196 8076 202
rect 7626 190 8024 196
rect 7626 -960 7738 190
rect 8024 138 8076 144
rect 8730 -960 8842 480
rect 9772 400 9824 406
rect 9926 354 10038 480
rect 9824 348 10038 354
rect 9772 342 10038 348
rect 9784 326 10038 342
rect 9926 -960 10038 326
rect 11122 -960 11234 480
rect 15948 480 15976 614
rect 17052 480 17080 682
rect 18052 536 18104 542
rect 12162 439 12218 448
rect 12176 354 12204 439
rect 12318 354 12430 480
rect 12176 326 12430 354
rect 12318 -960 12430 326
rect 13514 354 13626 480
rect 14556 468 14608 474
rect 14556 410 14608 416
rect 13726 368 13782 377
rect 13514 326 13726 354
rect 13514 -960 13626 326
rect 14568 354 14596 410
rect 14710 354 14822 480
rect 14568 326 14822 354
rect 13726 303 13782 312
rect 14710 -960 14822 326
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18052 478 18104 484
rect 19444 480 19472 886
rect 18064 354 18092 478
rect 18206 354 18318 480
rect 18064 326 18318 354
rect 18206 -960 18318 326
rect 19402 -960 19514 480
rect 19812 66 19840 3060
rect 20598 82 20710 480
rect 20916 134 20944 3060
rect 21824 876 21876 882
rect 21824 818 21876 824
rect 21836 480 21864 818
rect 20456 66 20710 82
rect 20904 128 20956 134
rect 20904 70 20956 76
rect 19800 60 19852 66
rect 19800 2 19852 8
rect 20444 60 20710 66
rect 20496 54 20710 60
rect 20444 2 20496 8
rect 20598 -960 20710 54
rect 21794 -960 21906 480
rect 22020 338 22048 3060
rect 22990 354 23102 480
rect 22848 338 23102 354
rect 22008 332 22060 338
rect 22008 274 22060 280
rect 22836 332 23102 338
rect 22888 326 23102 332
rect 22836 274 22888 280
rect 22990 -960 23102 326
rect 23216 270 23244 3060
rect 23952 3046 24242 3074
rect 25056 3046 25346 3074
rect 26344 3046 26450 3074
rect 23204 264 23256 270
rect 23204 206 23256 212
rect 23952 105 23980 3046
rect 24186 218 24298 480
rect 24584 264 24636 270
rect 24186 212 24584 218
rect 25056 241 25084 3046
rect 24186 206 24636 212
rect 25042 232 25098 241
rect 24186 190 24624 206
rect 23938 96 23994 105
rect 23938 31 23994 40
rect 24186 -960 24298 190
rect 25042 167 25098 176
rect 25290 218 25402 480
rect 25686 232 25742 241
rect 25290 190 25686 218
rect 25290 -960 25402 190
rect 26344 202 26372 3046
rect 26608 2984 26660 2990
rect 26608 2926 26660 2932
rect 26620 1578 26648 2926
rect 26528 1550 26648 1578
rect 26528 480 26556 1550
rect 27540 814 27568 3060
rect 27712 2916 27764 2922
rect 27712 2858 27764 2864
rect 27528 808 27580 814
rect 27528 750 27580 756
rect 27724 480 27752 2858
rect 25686 167 25742 176
rect 26332 196 26384 202
rect 26332 138 26384 144
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28644 406 28672 3060
rect 28906 640 28962 649
rect 29748 610 29776 3060
rect 28906 575 28962 584
rect 29736 604 29788 610
rect 28920 480 28948 575
rect 29736 546 29788 552
rect 30852 513 30880 3060
rect 30838 504 30894 513
rect 28632 400 28684 406
rect 28632 342 28684 348
rect 28878 -960 28990 480
rect 30074 218 30186 480
rect 30838 439 30894 448
rect 30074 202 30328 218
rect 30074 196 30340 202
rect 30074 190 30288 196
rect 30074 -960 30186 190
rect 30288 138 30340 144
rect 31116 128 31168 134
rect 31270 82 31382 480
rect 31956 377 31984 3060
rect 32220 400 32272 406
rect 31942 368 31998 377
rect 32374 354 32486 480
rect 33060 474 33088 3060
rect 33600 2848 33652 2854
rect 33600 2790 33652 2796
rect 33612 480 33640 2790
rect 34164 678 34192 3060
rect 35268 746 35296 3060
rect 35256 740 35308 746
rect 35256 682 35308 688
rect 34152 672 34204 678
rect 34152 614 34204 620
rect 35992 672 36044 678
rect 35992 614 36044 620
rect 36004 480 36032 614
rect 36372 542 36400 3060
rect 37476 950 37504 3060
rect 38212 3046 38594 3074
rect 37464 944 37516 950
rect 37464 886 37516 892
rect 36360 536 36412 542
rect 33048 468 33100 474
rect 33048 410 33100 416
rect 32272 348 32486 354
rect 32220 342 32486 348
rect 32232 326 32486 342
rect 31942 303 31998 312
rect 31168 76 31382 82
rect 31116 70 31382 76
rect 31128 54 31382 70
rect 31270 -960 31382 54
rect 32374 -960 32486 326
rect 33570 -960 33682 480
rect 34612 468 34664 474
rect 34612 410 34664 416
rect 34624 354 34652 410
rect 34766 354 34878 480
rect 34624 326 34878 354
rect 34766 -960 34878 326
rect 35962 -960 36074 480
rect 36360 478 36412 484
rect 37002 96 37058 105
rect 37158 82 37270 480
rect 37058 54 37270 82
rect 38212 66 38240 3046
rect 39684 882 39712 3060
rect 40512 3046 40802 3074
rect 40960 3062 41012 3068
rect 39672 876 39724 882
rect 39672 818 39724 824
rect 39580 604 39632 610
rect 39580 546 39632 552
rect 38568 536 38620 542
rect 38354 354 38466 480
rect 38568 478 38620 484
rect 39592 480 39620 546
rect 38580 354 38608 478
rect 38354 326 38608 354
rect 37002 31 37058 40
rect 37158 -960 37270 54
rect 38200 60 38252 66
rect 38200 2 38252 8
rect 38354 -960 38466 326
rect 39550 -960 39662 480
rect 40512 338 40540 3046
rect 40972 1578 41000 3062
rect 40696 1550 41000 1578
rect 41616 3046 41906 3074
rect 42812 3046 43010 3074
rect 40696 480 40724 1550
rect 40500 332 40552 338
rect 40500 274 40552 280
rect 40654 -960 40766 480
rect 41616 270 41644 3046
rect 41604 264 41656 270
rect 41604 206 41656 212
rect 41850 218 41962 480
rect 42248 264 42300 270
rect 41850 212 42248 218
rect 41850 206 42300 212
rect 42706 232 42762 241
rect 41850 190 42288 206
rect 41850 -960 41962 190
rect 42812 218 42840 3046
rect 44100 2990 44128 3060
rect 44088 2984 44140 2990
rect 44088 2926 44140 2932
rect 44272 2984 44324 2990
rect 44272 2926 44324 2932
rect 44284 480 44312 2926
rect 45204 2922 45232 3060
rect 45192 2916 45244 2922
rect 45192 2858 45244 2864
rect 46308 649 46336 3060
rect 46294 640 46350 649
rect 46294 575 46350 584
rect 43046 354 43158 480
rect 42904 338 43158 354
rect 42892 332 43158 338
rect 42944 326 43158 332
rect 42892 274 42944 280
rect 42762 190 42840 218
rect 42706 167 42762 176
rect 43046 -960 43158 326
rect 44242 -960 44354 480
rect 45438 82 45550 480
rect 45296 66 45550 82
rect 45284 60 45550 66
rect 45336 54 45550 60
rect 45284 2 45336 8
rect 45438 -960 45550 54
rect 46634 218 46746 480
rect 46846 232 46902 241
rect 46634 190 46846 218
rect 46634 -960 46746 190
rect 47412 202 47440 3060
rect 47860 2984 47912 2990
rect 47860 2926 47912 2932
rect 47872 480 47900 2926
rect 46846 167 46902 176
rect 47400 196 47452 202
rect 47400 138 47452 144
rect 47830 -960 47942 480
rect 48516 134 48544 3060
rect 48976 480 49004 3606
rect 51356 3460 51408 3466
rect 51356 3402 51408 3408
rect 48504 128 48556 134
rect 48504 70 48556 76
rect 48934 -960 49046 480
rect 49620 406 49648 3060
rect 50160 3052 50212 3058
rect 50160 2994 50212 3000
rect 50172 480 50200 2994
rect 50724 2854 50752 3060
rect 50712 2848 50764 2854
rect 50712 2790 50764 2796
rect 51368 480 51396 3402
rect 49608 400 49660 406
rect 49608 342 49660 348
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 51828 474 51856 3060
rect 52564 480 52592 3674
rect 54944 3528 54996 3534
rect 54944 3470 54996 3476
rect 52932 678 52960 3060
rect 52920 672 52972 678
rect 52920 614 52972 620
rect 51816 468 51868 474
rect 51816 410 51868 416
rect 52522 -960 52634 480
rect 53564 128 53616 134
rect 53718 82 53830 480
rect 54036 105 54064 3060
rect 54956 480 54984 3470
rect 55140 542 55168 3060
rect 55128 536 55180 542
rect 53616 76 53830 82
rect 53564 70 53830 76
rect 53576 54 53830 70
rect 53718 -960 53830 54
rect 54022 96 54078 105
rect 54022 31 54078 40
rect 54914 -960 55026 480
rect 55128 478 55180 484
rect 56060 480 56088 3742
rect 64788 3664 64840 3670
rect 64840 3612 65090 3618
rect 64788 3606 65090 3612
rect 60832 3596 60884 3602
rect 64800 3590 65090 3606
rect 60832 3538 60884 3544
rect 58808 3256 58860 3262
rect 58808 3198 58860 3204
rect 56968 3188 57020 3194
rect 56968 3130 57020 3136
rect 56244 610 56272 3060
rect 56232 604 56284 610
rect 56232 546 56284 552
rect 56018 -960 56130 480
rect 56980 354 57008 3130
rect 57060 3120 57112 3126
rect 57112 3068 57362 3074
rect 57060 3062 57362 3068
rect 57072 3046 57362 3062
rect 58176 3046 58466 3074
rect 57214 354 57326 480
rect 56980 326 57326 354
rect 57214 -960 57326 326
rect 58176 270 58204 3046
rect 58410 354 58522 480
rect 58820 354 58848 3198
rect 58410 326 58848 354
rect 59372 3046 59570 3074
rect 59372 338 59400 3046
rect 60660 2922 60688 3060
rect 60648 2916 60700 2922
rect 60648 2858 60700 2864
rect 59636 2848 59688 2854
rect 59636 2790 59688 2796
rect 59648 480 59676 2790
rect 60844 480 60872 3538
rect 63224 3392 63276 3398
rect 63224 3334 63276 3340
rect 62028 3324 62080 3330
rect 62028 3266 62080 3272
rect 59360 332 59412 338
rect 58164 264 58216 270
rect 58164 206 58216 212
rect 58410 -960 58522 326
rect 59360 274 59412 280
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61764 66 61792 3060
rect 62040 480 62068 3266
rect 61752 60 61804 66
rect 61752 2 61804 8
rect 61998 -960 62110 480
rect 62868 241 62896 3060
rect 63236 480 63264 3334
rect 63420 3046 63986 3074
rect 63420 2990 63448 3046
rect 63408 2984 63460 2990
rect 63408 2926 63460 2932
rect 64328 2848 64380 2854
rect 64328 2790 64380 2796
rect 64340 480 64368 2790
rect 65536 480 65564 3810
rect 71412 3800 71464 3806
rect 68112 3738 68402 3754
rect 90088 3800 90140 3806
rect 71464 3748 71714 3754
rect 71412 3742 71714 3748
rect 68100 3732 68402 3738
rect 68152 3726 68402 3732
rect 71424 3726 71714 3742
rect 85776 3738 86066 3754
rect 90088 3742 90140 3748
rect 71872 3732 71924 3738
rect 68100 3674 68152 3680
rect 71872 3674 71924 3680
rect 85764 3732 86066 3738
rect 85816 3726 86066 3732
rect 86868 3732 86920 3738
rect 85764 3674 85816 3680
rect 86868 3674 86920 3680
rect 66720 3664 66772 3670
rect 66720 3606 66772 3612
rect 65904 3058 66194 3074
rect 65892 3052 66194 3058
rect 65944 3046 66194 3052
rect 65892 2994 65944 3000
rect 66732 480 66760 3606
rect 71884 3534 71912 3674
rect 81440 3664 81492 3670
rect 75932 3602 76130 3618
rect 84476 3664 84528 3670
rect 81492 3612 81650 3618
rect 81440 3606 81650 3612
rect 84476 3606 84528 3612
rect 75920 3596 76130 3602
rect 75972 3590 76130 3596
rect 76288 3596 76340 3602
rect 75920 3538 75972 3544
rect 81452 3590 81650 3606
rect 76288 3538 76340 3544
rect 70308 3528 70360 3534
rect 67008 3466 67298 3482
rect 71504 3528 71556 3534
rect 70360 3476 70610 3482
rect 70308 3470 70610 3476
rect 71504 3470 71556 3476
rect 71872 3528 71924 3534
rect 71872 3470 71924 3476
rect 72976 3528 73028 3534
rect 72976 3470 73028 3476
rect 66996 3460 67298 3466
rect 67048 3454 67298 3460
rect 70124 3460 70176 3466
rect 66996 3402 67048 3408
rect 70320 3454 70610 3470
rect 70124 3402 70176 3408
rect 69112 3052 69164 3058
rect 69112 2994 69164 3000
rect 67916 2984 67968 2990
rect 67916 2926 67968 2932
rect 67928 480 67956 2926
rect 68836 2848 68888 2854
rect 68836 2790 68888 2796
rect 68848 1222 68876 2790
rect 68836 1216 68888 1222
rect 68836 1158 68888 1164
rect 69124 480 69152 2994
rect 62854 232 62910 241
rect 62854 167 62910 176
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 69492 134 69520 3060
rect 70136 218 70164 3402
rect 71516 480 71544 3470
rect 72528 3194 72818 3210
rect 72516 3188 72818 3194
rect 72568 3182 72818 3188
rect 72516 3130 72568 3136
rect 70278 218 70390 480
rect 70136 190 70390 218
rect 69480 128 69532 134
rect 69480 70 69532 76
rect 70278 -960 70390 190
rect 71474 -960 71586 480
rect 72578 354 72690 480
rect 72988 354 73016 3470
rect 73632 3318 73922 3346
rect 73632 3262 73660 3318
rect 73620 3256 73672 3262
rect 73620 3198 73672 3204
rect 73804 3188 73856 3194
rect 73804 3130 73856 3136
rect 73816 480 73844 3130
rect 75012 2922 75040 3060
rect 75000 2916 75052 2922
rect 75000 2858 75052 2864
rect 75368 2916 75420 2922
rect 75368 2858 75420 2864
rect 72578 326 73016 354
rect 72578 -960 72690 326
rect 73774 -960 73886 480
rect 74970 354 75082 480
rect 75380 354 75408 2858
rect 76300 1850 76328 3538
rect 78036 3392 78088 3398
rect 76944 3330 77234 3346
rect 83280 3392 83332 3398
rect 78088 3340 78338 3346
rect 78036 3334 78338 3340
rect 83280 3334 83332 3340
rect 76932 3324 77234 3330
rect 76984 3318 77234 3324
rect 78048 3318 78338 3334
rect 82084 3324 82136 3330
rect 76932 3266 76984 3272
rect 82084 3266 82136 3272
rect 77392 3256 77444 3262
rect 77392 3198 77444 3204
rect 77116 2984 77168 2990
rect 77116 2926 77168 2932
rect 76208 1822 76328 1850
rect 76208 480 76236 1822
rect 77128 1358 77156 2926
rect 77116 1352 77168 1358
rect 77116 1294 77168 1300
rect 77404 480 77432 3198
rect 80888 3120 80940 3126
rect 80888 3062 80940 3068
rect 78588 2984 78640 2990
rect 78588 2926 78640 2932
rect 78600 480 78628 2926
rect 79428 1222 79456 3060
rect 79692 2848 79744 2854
rect 79692 2790 79744 2796
rect 79416 1216 79468 1222
rect 79416 1158 79468 1164
rect 79704 480 79732 2790
rect 80900 480 80928 3062
rect 82096 480 82124 3266
rect 82740 1358 82768 3060
rect 82728 1352 82780 1358
rect 82728 1294 82780 1300
rect 83292 480 83320 3334
rect 83568 3058 83858 3074
rect 83556 3052 83858 3058
rect 83608 3046 83858 3052
rect 83556 2994 83608 3000
rect 84488 480 84516 3606
rect 84672 3466 84962 3482
rect 84660 3460 84962 3466
rect 84712 3454 84962 3460
rect 84660 3402 84712 3408
rect 85488 2916 85540 2922
rect 85488 2858 85540 2864
rect 85672 2916 85724 2922
rect 85672 2858 85724 2864
rect 85500 1290 85528 2858
rect 85488 1284 85540 1290
rect 85488 1226 85540 1232
rect 85684 480 85712 2858
rect 86880 480 86908 3674
rect 86960 3528 87012 3534
rect 87788 3528 87840 3534
rect 87012 3476 87170 3482
rect 86960 3470 87170 3476
rect 87788 3470 87840 3476
rect 86972 3454 87170 3470
rect 74970 326 75408 354
rect 74970 -960 75082 326
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87800 218 87828 3470
rect 89536 3460 89588 3466
rect 89536 3402 89588 3408
rect 87984 3194 88274 3210
rect 87972 3188 88274 3194
rect 88024 3182 88274 3188
rect 87972 3130 88024 3136
rect 88984 2984 89036 2990
rect 88984 2926 89036 2932
rect 88996 1358 89024 2926
rect 88984 1352 89036 1358
rect 88984 1294 89036 1300
rect 89364 1290 89392 3060
rect 89352 1284 89404 1290
rect 89352 1226 89404 1232
rect 87942 218 88054 480
rect 87800 190 88054 218
rect 87942 -960 88054 190
rect 89138 354 89250 480
rect 89548 354 89576 3402
rect 89138 326 89576 354
rect 90100 354 90128 3742
rect 90192 3602 90482 3618
rect 97644 3602 97672 3810
rect 103428 3800 103480 3806
rect 100128 3738 100418 3754
rect 104348 3800 104400 3806
rect 103480 3748 103730 3754
rect 103428 3742 103730 3748
rect 104348 3742 104400 3748
rect 100116 3732 100418 3738
rect 100168 3726 100418 3732
rect 103440 3726 103730 3742
rect 100116 3674 100168 3680
rect 97908 3664 97960 3670
rect 97960 3612 98210 3618
rect 97908 3606 98210 3612
rect 90180 3596 90482 3602
rect 90232 3590 90482 3596
rect 97632 3596 97684 3602
rect 90180 3538 90232 3544
rect 97920 3590 98210 3606
rect 97632 3538 97684 3544
rect 97448 3528 97500 3534
rect 97448 3470 97500 3476
rect 98644 3528 98696 3534
rect 98644 3470 98696 3476
rect 92940 3392 92992 3398
rect 92940 3334 92992 3340
rect 93952 3392 94004 3398
rect 93952 3334 94004 3340
rect 91284 3256 91336 3262
rect 91336 3204 91586 3210
rect 91284 3198 91586 3204
rect 91296 3182 91586 3198
rect 92848 3188 92900 3194
rect 92848 3130 92900 3136
rect 92400 3058 92690 3074
rect 92388 3052 92690 3058
rect 92440 3046 92690 3052
rect 92388 2994 92440 3000
rect 91928 2848 91980 2854
rect 91928 2790 91980 2796
rect 90334 354 90446 480
rect 90100 326 90446 354
rect 89138 -960 89250 326
rect 90334 -960 90446 326
rect 91530 354 91642 480
rect 91940 354 91968 2790
rect 92860 1578 92888 3130
rect 92768 1550 92888 1578
rect 92768 480 92796 1550
rect 92952 1290 92980 3334
rect 93780 1358 93808 3060
rect 93768 1352 93820 1358
rect 93768 1294 93820 1300
rect 92940 1284 92992 1290
rect 92940 1226 92992 1232
rect 93964 480 93992 3334
rect 95712 3330 96002 3346
rect 95700 3324 96002 3330
rect 95752 3318 96002 3324
rect 95700 3266 95752 3272
rect 96252 3256 96304 3262
rect 96252 3198 96304 3204
rect 94596 3120 94648 3126
rect 94648 3068 94898 3074
rect 94596 3062 94898 3068
rect 94608 3046 94898 3062
rect 95148 3052 95200 3058
rect 95148 2994 95200 3000
rect 95056 2916 95108 2922
rect 95056 2858 95108 2864
rect 95068 1204 95096 2858
rect 95160 1358 95188 2994
rect 95148 1352 95200 1358
rect 95148 1294 95200 1300
rect 95068 1176 95188 1204
rect 95160 480 95188 1176
rect 96264 480 96292 3198
rect 97092 1290 97120 3060
rect 97080 1284 97132 1290
rect 97080 1226 97132 1232
rect 97460 480 97488 3470
rect 98656 480 98684 3470
rect 102336 3466 102626 3482
rect 102324 3460 102626 3466
rect 102376 3454 102626 3460
rect 102324 3402 102376 3408
rect 101036 3392 101088 3398
rect 101036 3334 101088 3340
rect 99300 1358 99328 3060
rect 99840 2848 99892 2854
rect 99840 2790 99892 2796
rect 99288 1352 99340 1358
rect 99288 1294 99340 1300
rect 99852 480 99880 2790
rect 101048 480 101076 3334
rect 103336 3324 103388 3330
rect 103336 3266 103388 3272
rect 102232 2984 102284 2990
rect 102232 2926 102284 2932
rect 102244 480 102272 2926
rect 103348 480 103376 3266
rect 91530 326 91968 354
rect 91530 -960 91642 326
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104360 218 104388 3742
rect 116688 3738 116978 3754
rect 106648 3732 106700 3738
rect 106648 3674 106700 3680
rect 116676 3732 116978 3738
rect 116728 3726 116978 3732
rect 116676 3674 116728 3680
rect 105636 3120 105688 3126
rect 104544 3058 104834 3074
rect 106096 3120 106148 3126
rect 105688 3068 105938 3074
rect 105636 3062 105938 3068
rect 106096 3062 106148 3068
rect 104532 3052 104834 3058
rect 104584 3046 104834 3052
rect 105648 3046 105938 3062
rect 104532 2994 104584 3000
rect 104502 218 104614 480
rect 104360 190 104614 218
rect 104502 -960 104614 190
rect 105698 354 105810 480
rect 106108 354 106136 3062
rect 105698 326 106136 354
rect 106660 354 106688 3674
rect 110052 3664 110104 3670
rect 118884 3664 118936 3670
rect 110104 3612 110354 3618
rect 110052 3606 110354 3612
rect 125968 3664 126020 3670
rect 118936 3612 119186 3618
rect 118884 3606 119186 3612
rect 108488 3596 108540 3602
rect 110064 3590 110354 3606
rect 118896 3590 119186 3606
rect 120000 3602 120290 3618
rect 136548 3664 136600 3670
rect 125968 3606 126020 3612
rect 119988 3596 120290 3602
rect 108488 3538 108540 3544
rect 120040 3590 120290 3596
rect 122288 3596 122340 3602
rect 119988 3538 120040 3544
rect 122288 3538 122340 3544
rect 106740 3256 106792 3262
rect 106792 3204 107042 3210
rect 106740 3198 107042 3204
rect 106752 3182 107042 3198
rect 107856 3046 108146 3074
rect 107856 2922 107884 3046
rect 107844 2916 107896 2922
rect 107844 2858 107896 2864
rect 106894 354 107006 480
rect 106660 326 107006 354
rect 105698 -960 105810 326
rect 106894 -960 107006 326
rect 108090 354 108202 480
rect 108500 354 108528 3538
rect 110512 3528 110564 3534
rect 110512 3470 110564 3476
rect 108960 3194 109250 3210
rect 108948 3188 109250 3194
rect 109000 3182 109250 3188
rect 109408 3188 109460 3194
rect 108948 3130 109000 3136
rect 109408 3130 109460 3136
rect 109420 1578 109448 3130
rect 109328 1550 109448 1578
rect 109328 480 109356 1550
rect 110524 480 110552 3470
rect 111168 3466 111458 3482
rect 111156 3460 111458 3466
rect 111208 3454 111458 3460
rect 117596 3460 117648 3466
rect 111156 3402 111208 3408
rect 117596 3402 117648 3408
rect 113364 3392 113416 3398
rect 116400 3392 116452 3398
rect 113416 3340 113666 3346
rect 113364 3334 113666 3340
rect 113376 3318 113666 3334
rect 115584 3330 115874 3346
rect 116400 3334 116452 3340
rect 115572 3324 115874 3330
rect 115624 3318 115874 3324
rect 115572 3266 115624 3272
rect 111616 3256 111668 3262
rect 111616 3198 111668 3204
rect 111628 480 111656 3198
rect 112272 3046 112562 3074
rect 112812 3052 112864 3058
rect 112272 2854 112300 3046
rect 112812 2994 112864 3000
rect 114572 3046 114770 3074
rect 112260 2848 112312 2854
rect 112260 2790 112312 2796
rect 112824 480 112852 2994
rect 114008 2984 114060 2990
rect 114008 2926 114060 2932
rect 114020 480 114048 2926
rect 114572 2922 114600 3046
rect 114560 2916 114612 2922
rect 114560 2858 114612 2864
rect 115204 2916 115256 2922
rect 115204 2858 115256 2864
rect 115216 480 115244 2858
rect 116412 480 116440 3334
rect 117608 480 117636 3402
rect 121552 3392 121604 3398
rect 121552 3334 121604 3340
rect 119896 3324 119948 3330
rect 119896 3266 119948 3272
rect 117780 3120 117832 3126
rect 117832 3068 118082 3074
rect 117780 3062 118082 3068
rect 117792 3046 118082 3062
rect 118792 2848 118844 2854
rect 118792 2790 118844 2796
rect 118804 480 118832 2790
rect 119908 480 119936 3266
rect 121104 3194 121394 3210
rect 121092 3188 121394 3194
rect 121144 3182 121394 3188
rect 121092 3130 121144 3136
rect 121564 3126 121592 3334
rect 121184 3120 121236 3126
rect 121184 3062 121236 3068
rect 121552 3120 121604 3126
rect 121552 3062 121604 3068
rect 121196 1578 121224 3062
rect 121104 1550 121224 1578
rect 121104 480 121132 1550
rect 122300 480 122328 3538
rect 122380 3528 122432 3534
rect 122432 3476 122498 3482
rect 122380 3470 122498 3476
rect 122392 3454 122498 3470
rect 123300 3256 123352 3262
rect 123760 3256 123812 3262
rect 123352 3204 123602 3210
rect 123300 3198 123602 3204
rect 123760 3198 123812 3204
rect 123312 3182 123602 3198
rect 123772 1714 123800 3198
rect 124416 3058 124706 3074
rect 124404 3052 124706 3058
rect 124456 3046 124706 3052
rect 125048 3052 125100 3058
rect 124404 2994 124456 3000
rect 125048 2994 125100 3000
rect 125612 3046 125810 3074
rect 123496 1686 123800 1714
rect 123496 480 123524 1686
rect 108090 326 108528 354
rect 108090 -960 108202 326
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 354 124762 480
rect 125060 354 125088 2994
rect 125612 2990 125640 3046
rect 125600 2984 125652 2990
rect 125600 2926 125652 2932
rect 125980 1850 126008 3606
rect 133248 3602 133538 3618
rect 143632 3664 143684 3670
rect 136600 3612 136850 3618
rect 136548 3606 136850 3612
rect 153200 3664 153252 3670
rect 143632 3606 143684 3612
rect 133236 3596 133538 3602
rect 133288 3590 133538 3596
rect 136560 3590 136850 3606
rect 142528 3596 142580 3602
rect 133236 3538 133288 3544
rect 142528 3538 142580 3544
rect 129372 3528 129424 3534
rect 128832 3466 129122 3482
rect 139860 3528 139912 3534
rect 129372 3470 129424 3476
rect 128820 3460 129122 3466
rect 128872 3454 129122 3460
rect 128820 3402 128872 3408
rect 128176 3392 128228 3398
rect 128176 3334 128228 3340
rect 127716 3120 127768 3126
rect 126624 3046 126914 3074
rect 127768 3068 128018 3074
rect 127716 3062 128018 3068
rect 127728 3046 128018 3062
rect 126624 2922 126652 3046
rect 126612 2916 126664 2922
rect 126612 2858 126664 2864
rect 126980 2916 127032 2922
rect 126980 2858 127032 2864
rect 125888 1822 126008 1850
rect 125888 480 125916 1822
rect 126992 480 127020 2858
rect 128188 480 128216 3334
rect 129384 480 129412 3470
rect 138768 3466 139058 3482
rect 141608 3528 141660 3534
rect 139912 3476 140162 3482
rect 139860 3470 140162 3476
rect 141608 3470 141660 3476
rect 138756 3460 139058 3466
rect 138808 3454 139058 3460
rect 139872 3454 140162 3470
rect 138756 3402 138808 3408
rect 130568 3392 130620 3398
rect 140688 3392 140740 3398
rect 130568 3334 130620 3340
rect 129660 3046 130226 3074
rect 129660 2854 129688 3046
rect 129648 2848 129700 2854
rect 129648 2790 129700 2796
rect 130580 480 130608 3334
rect 131040 3330 131330 3346
rect 140740 3340 141266 3346
rect 140688 3334 141266 3340
rect 131028 3324 131330 3330
rect 131080 3318 131330 3324
rect 140044 3324 140096 3330
rect 131028 3266 131080 3272
rect 140700 3318 141266 3334
rect 140044 3266 140096 3272
rect 134340 3256 134392 3262
rect 132144 3194 132434 3210
rect 137652 3256 137704 3262
rect 134392 3204 134642 3210
rect 134340 3198 134642 3204
rect 137652 3198 137704 3204
rect 132132 3188 132434 3194
rect 132184 3182 132434 3188
rect 134352 3182 134642 3198
rect 136456 3188 136508 3194
rect 132132 3130 132184 3136
rect 136456 3130 136508 3136
rect 131764 3120 131816 3126
rect 131764 3062 131816 3068
rect 131776 480 131804 3062
rect 135180 3058 135746 3074
rect 135168 3052 135746 3058
rect 135220 3046 135746 3052
rect 135904 3052 135956 3058
rect 135168 2994 135220 3000
rect 135904 2994 135956 3000
rect 134156 2984 134208 2990
rect 134156 2926 134208 2932
rect 132960 2848 133012 2854
rect 132960 2790 133012 2796
rect 132972 480 133000 2790
rect 134168 480 134196 2926
rect 135916 1578 135944 2994
rect 135272 1550 135944 1578
rect 135272 480 135300 1550
rect 136468 480 136496 3130
rect 137664 480 137692 3198
rect 137940 2922 137968 3060
rect 137928 2916 137980 2922
rect 137928 2858 137980 2864
rect 138848 2916 138900 2922
rect 138848 2858 138900 2864
rect 138860 480 138888 2858
rect 140056 480 140084 3266
rect 124650 326 125088 354
rect 124650 -960 124762 326
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 354 141322 480
rect 141620 354 141648 3470
rect 142068 3120 142120 3126
rect 142120 3068 142370 3074
rect 142068 3062 142370 3068
rect 142080 3046 142370 3062
rect 142540 1850 142568 3538
rect 143460 2854 143488 3060
rect 143448 2848 143500 2854
rect 143448 2790 143500 2796
rect 143644 1850 143672 3606
rect 152016 3602 152306 3618
rect 153252 3612 153410 3618
rect 153200 3606 153410 3612
rect 152004 3596 152306 3602
rect 152056 3590 152306 3596
rect 153212 3590 153410 3606
rect 152004 3538 152056 3544
rect 150900 3528 150952 3534
rect 149808 3466 150098 3482
rect 150952 3476 151202 3482
rect 150900 3470 151202 3476
rect 149796 3460 150098 3466
rect 149848 3454 150098 3460
rect 150912 3454 151202 3470
rect 149796 3402 149848 3408
rect 147588 3392 147640 3398
rect 154028 3392 154080 3398
rect 147640 3340 147890 3346
rect 147588 3334 147890 3340
rect 163044 3392 163096 3398
rect 154028 3334 154080 3340
rect 145932 3324 145984 3330
rect 147600 3318 147890 3334
rect 145932 3266 145984 3272
rect 144736 3120 144788 3126
rect 144736 3062 144788 3068
rect 144564 2990 144592 3060
rect 144552 2984 144604 2990
rect 144552 2926 144604 2932
rect 142448 1822 142568 1850
rect 143552 1822 143672 1850
rect 142448 480 142476 1822
rect 143552 480 143580 1822
rect 144748 480 144776 3062
rect 145392 3058 145682 3074
rect 145380 3052 145682 3058
rect 145432 3046 145682 3052
rect 145380 2994 145432 3000
rect 145944 480 145972 3266
rect 151820 3256 151872 3262
rect 146220 3194 146786 3210
rect 151820 3198 151872 3204
rect 146208 3188 146786 3194
rect 146260 3182 146786 3188
rect 146208 3130 146260 3136
rect 149520 3120 149572 3126
rect 149520 3062 149572 3068
rect 147128 3052 147180 3058
rect 147128 2994 147180 3000
rect 147140 480 147168 2994
rect 148980 2990 149008 3060
rect 148968 2984 149020 2990
rect 148968 2926 149020 2932
rect 148324 2916 148376 2922
rect 148324 2858 148376 2864
rect 148336 480 148364 2858
rect 149532 480 149560 3062
rect 150624 2848 150676 2854
rect 150624 2790 150676 2796
rect 150636 480 150664 2790
rect 151832 480 151860 3198
rect 153016 2984 153068 2990
rect 153016 2926 153068 2932
rect 153028 480 153056 2926
rect 141210 326 141648 354
rect 141210 -960 141322 326
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154040 218 154068 3334
rect 155328 3330 155618 3346
rect 166080 3392 166132 3398
rect 163096 3340 163346 3346
rect 163044 3334 163346 3340
rect 155316 3324 155618 3330
rect 155368 3318 155618 3324
rect 155776 3324 155828 3330
rect 155316 3266 155368 3272
rect 163056 3318 163346 3334
rect 164252 3330 164450 3346
rect 174084 3392 174136 3398
rect 166080 3334 166132 3340
rect 164240 3324 164450 3330
rect 155776 3266 155828 3272
rect 164292 3318 164450 3324
rect 164884 3324 164936 3330
rect 164240 3266 164292 3272
rect 164884 3266 164936 3272
rect 154224 3194 154514 3210
rect 154212 3188 154514 3194
rect 154264 3182 154514 3188
rect 154212 3130 154264 3136
rect 154182 218 154294 480
rect 154040 190 154294 218
rect 154182 -960 154294 190
rect 155378 354 155490 480
rect 155788 354 155816 3266
rect 160836 3256 160888 3262
rect 162492 3256 162544 3262
rect 160888 3204 161138 3210
rect 160836 3198 161138 3204
rect 162492 3198 162544 3204
rect 156328 3188 156380 3194
rect 160848 3182 161138 3198
rect 156328 3130 156380 3136
rect 155378 326 155816 354
rect 156340 354 156368 3130
rect 158720 3120 158772 3126
rect 156432 3058 156722 3074
rect 156420 3052 156722 3058
rect 156472 3046 156722 3052
rect 157536 3046 157826 3074
rect 160192 3120 160244 3126
rect 158772 3068 158930 3074
rect 158720 3062 158930 3068
rect 160192 3062 160244 3068
rect 158732 3046 158930 3062
rect 159272 3052 159324 3058
rect 156420 2994 156472 3000
rect 157536 2922 157564 3046
rect 159272 2994 159324 3000
rect 157524 2916 157576 2922
rect 157524 2858 157576 2864
rect 157800 2916 157852 2922
rect 157800 2858 157852 2864
rect 157812 480 157840 2858
rect 156574 354 156686 480
rect 156340 326 156686 354
rect 155378 -960 155490 326
rect 156574 -960 156686 326
rect 157770 -960 157882 480
rect 158874 354 158986 480
rect 159284 354 159312 2994
rect 160020 2854 160048 3060
rect 160008 2848 160060 2854
rect 160008 2790 160060 2796
rect 160204 1578 160232 3062
rect 162228 2990 162256 3060
rect 162216 2984 162268 2990
rect 162216 2926 162268 2932
rect 161296 2848 161348 2854
rect 161296 2790 161348 2796
rect 160112 1550 160232 1578
rect 160112 480 160140 1550
rect 161308 480 161336 2790
rect 162504 480 162532 3198
rect 163688 2984 163740 2990
rect 163688 2926 163740 2932
rect 163700 480 163728 2926
rect 164896 480 164924 3266
rect 165264 3194 165554 3210
rect 165252 3188 165554 3194
rect 165304 3182 165554 3188
rect 165712 3188 165764 3194
rect 165252 3130 165304 3136
rect 165712 3130 165764 3136
rect 165724 2990 165752 3130
rect 165712 2984 165764 2990
rect 165712 2926 165764 2932
rect 166092 480 166120 3334
rect 172992 3330 173282 3346
rect 183744 3392 183796 3398
rect 174136 3340 174386 3346
rect 174084 3334 174386 3340
rect 190644 3392 190696 3398
rect 183744 3334 183796 3340
rect 172980 3324 173282 3330
rect 173032 3318 173282 3324
rect 174096 3318 174386 3334
rect 176752 3324 176804 3330
rect 172980 3266 173032 3272
rect 176752 3266 176804 3272
rect 170772 3256 170824 3262
rect 171876 3256 171928 3262
rect 170824 3204 171074 3210
rect 170772 3198 171074 3204
rect 173164 3256 173216 3262
rect 171928 3204 172178 3210
rect 171876 3198 172178 3204
rect 173164 3198 173216 3204
rect 170784 3182 171074 3198
rect 171888 3182 172178 3198
rect 168564 3120 168616 3126
rect 166644 2922 166672 3060
rect 167472 3058 167762 3074
rect 168616 3068 168866 3074
rect 168564 3062 168866 3068
rect 167460 3052 167762 3058
rect 167512 3046 167762 3052
rect 168380 3052 168432 3058
rect 167460 2994 167512 3000
rect 168576 3046 168866 3062
rect 168380 2994 168432 3000
rect 167184 2984 167236 2990
rect 167184 2926 167236 2932
rect 166632 2916 166684 2922
rect 166632 2858 166684 2864
rect 167196 480 167224 2926
rect 168392 480 168420 2994
rect 169576 2916 169628 2922
rect 169576 2858 169628 2864
rect 169588 480 169616 2858
rect 169956 2854 169984 3060
rect 171968 2984 172020 2990
rect 171968 2926 172020 2932
rect 169944 2848 169996 2854
rect 169944 2790 169996 2796
rect 170772 2848 170824 2854
rect 170772 2790 170824 2796
rect 170784 480 170812 2790
rect 171980 480 172008 2926
rect 173176 480 173204 3198
rect 174268 3188 174320 3194
rect 174268 3130 174320 3136
rect 174280 480 174308 3130
rect 176292 3120 176344 3126
rect 175292 3058 175490 3074
rect 176344 3068 176594 3074
rect 176292 3062 176594 3068
rect 175280 3052 175490 3058
rect 175332 3046 175490 3052
rect 175832 3052 175884 3058
rect 175280 2994 175332 3000
rect 176304 3046 176594 3062
rect 175832 2994 175884 3000
rect 158874 326 159312 354
rect 158874 -960 158986 326
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 354 175546 480
rect 175844 354 175872 2994
rect 176764 1714 176792 3266
rect 180892 3256 180944 3262
rect 181444 3256 181496 3262
rect 180944 3204 181010 3210
rect 180892 3198 181010 3204
rect 181444 3198 181496 3204
rect 179052 3188 179104 3194
rect 180904 3182 181010 3198
rect 179052 3130 179104 3136
rect 177684 2922 177712 3060
rect 177672 2916 177724 2922
rect 177672 2858 177724 2864
rect 177856 2916 177908 2922
rect 177856 2858 177908 2864
rect 176672 1686 176792 1714
rect 176672 480 176700 1686
rect 177868 480 177896 2858
rect 178788 2854 178816 3060
rect 178776 2848 178828 2854
rect 178776 2790 178828 2796
rect 179064 480 179092 3130
rect 179892 2990 179920 3060
rect 179880 2984 179932 2990
rect 179880 2926 179932 2932
rect 180248 2848 180300 2854
rect 180248 2790 180300 2796
rect 180260 480 180288 2790
rect 181456 480 181484 3198
rect 181812 3120 181864 3126
rect 181864 3068 182114 3074
rect 181812 3062 182114 3068
rect 181824 3046 182114 3062
rect 182928 3058 183218 3074
rect 182916 3052 183218 3058
rect 182968 3046 183218 3052
rect 182916 2994 182968 3000
rect 182548 2984 182600 2990
rect 182548 2926 182600 2932
rect 182560 480 182588 2926
rect 183756 480 183784 3334
rect 184032 3330 184322 3346
rect 553308 3392 553360 3398
rect 190696 3340 190946 3346
rect 190644 3334 190946 3340
rect 184020 3324 184322 3330
rect 184072 3318 184322 3324
rect 184940 3324 184992 3330
rect 184020 3266 184072 3272
rect 190656 3318 190946 3334
rect 549838 3330 550128 3346
rect 553150 3340 553308 3346
rect 553150 3334 553360 3340
rect 571524 3392 571576 3398
rect 571524 3334 571576 3340
rect 549838 3324 550140 3330
rect 549838 3318 550088 3324
rect 184940 3266 184992 3272
rect 553150 3318 553348 3334
rect 568028 3324 568080 3330
rect 550088 3266 550140 3272
rect 568028 3266 568080 3272
rect 184952 480 184980 3266
rect 188436 3256 188488 3262
rect 186332 3194 186530 3210
rect 191840 3256 191892 3262
rect 188488 3204 188738 3210
rect 188436 3198 188738 3204
rect 197360 3256 197412 3262
rect 191892 3204 192050 3210
rect 191840 3198 192050 3204
rect 214472 3256 214524 3262
rect 197412 3204 197570 3210
rect 197360 3198 197570 3204
rect 186320 3188 186530 3194
rect 186372 3182 186530 3188
rect 188448 3182 188738 3198
rect 190828 3188 190880 3194
rect 186320 3130 186372 3136
rect 191852 3182 192050 3198
rect 196808 3188 196860 3194
rect 190828 3130 190880 3136
rect 197372 3182 197570 3198
rect 202892 3194 203090 3210
rect 202880 3188 203090 3194
rect 196808 3130 196860 3136
rect 202932 3182 203090 3188
rect 206112 3182 206402 3210
rect 219348 3256 219400 3262
rect 214472 3198 214524 3204
rect 209872 3188 209924 3194
rect 202880 3130 202932 3136
rect 186136 3120 186188 3126
rect 186136 3062 186188 3068
rect 185412 2922 185440 3060
rect 185400 2916 185452 2922
rect 185400 2858 185452 2864
rect 186148 480 186176 3062
rect 187620 2922 187648 3060
rect 188528 3052 188580 3058
rect 188528 2994 188580 3000
rect 189552 3046 189842 3074
rect 187608 2916 187660 2922
rect 187608 2858 187660 2864
rect 187332 2848 187384 2854
rect 187332 2790 187384 2796
rect 187344 480 187372 2790
rect 188540 480 188568 2994
rect 189552 2990 189580 3046
rect 189540 2984 189592 2990
rect 189540 2926 189592 2932
rect 189724 2984 189776 2990
rect 189724 2926 189776 2932
rect 189736 480 189764 2926
rect 190840 480 190868 3130
rect 192852 3120 192904 3126
rect 193312 3120 193364 3126
rect 192904 3068 193154 3074
rect 192852 3062 193154 3068
rect 193312 3062 193364 3068
rect 192864 3046 193154 3062
rect 192392 2916 192444 2922
rect 192392 2858 192444 2864
rect 175434 326 175872 354
rect 175434 -960 175546 326
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 354 192106 480
rect 192404 354 192432 2858
rect 193324 1578 193352 3062
rect 194244 2854 194272 3060
rect 195072 3058 195362 3074
rect 195060 3052 195362 3058
rect 195112 3046 195362 3052
rect 195612 3052 195664 3058
rect 195060 2994 195112 3000
rect 195612 2994 195664 3000
rect 194232 2848 194284 2854
rect 194232 2790 194284 2796
rect 194416 2848 194468 2854
rect 194416 2790 194468 2796
rect 193232 1550 193352 1578
rect 193232 480 193260 1550
rect 194428 480 194456 2790
rect 195624 480 195652 2994
rect 196452 2990 196480 3060
rect 196440 2984 196492 2990
rect 196440 2926 196492 2932
rect 196820 480 196848 3130
rect 206112 3126 206140 3182
rect 209872 3130 209924 3136
rect 199476 3120 199528 3126
rect 198384 3046 198674 3074
rect 200304 3120 200356 3126
rect 199528 3068 199778 3074
rect 199476 3062 199778 3068
rect 206100 3120 206152 3126
rect 200304 3062 200356 3068
rect 199488 3046 199778 3062
rect 198384 2922 198412 3046
rect 198372 2916 198424 2922
rect 198372 2858 198424 2864
rect 199108 2916 199160 2922
rect 199108 2858 199160 2864
rect 198280 1352 198332 1358
rect 198280 1294 198332 1300
rect 191994 326 192432 354
rect 191994 -960 192106 326
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 354 197994 480
rect 198292 354 198320 1294
rect 199120 480 199148 2858
rect 200316 480 200344 3062
rect 200868 2854 200896 3060
rect 201696 3058 201986 3074
rect 201684 3052 201986 3058
rect 201736 3046 201986 3052
rect 201684 2994 201736 3000
rect 201500 2984 201552 2990
rect 201500 2926 201552 2932
rect 203892 2984 203944 2990
rect 203892 2926 203944 2932
rect 200856 2848 200908 2854
rect 200856 2790 200908 2796
rect 201512 480 201540 2926
rect 202696 2848 202748 2854
rect 202696 2790 202748 2796
rect 202708 480 202736 2790
rect 203904 480 203932 2926
rect 204180 1358 204208 3060
rect 205008 3046 205298 3074
rect 206100 3062 206152 3068
rect 206192 3120 206244 3126
rect 206192 3062 206244 3068
rect 205008 2922 205036 3046
rect 204996 2916 205048 2922
rect 204996 2858 205048 2864
rect 205088 2916 205140 2922
rect 205088 2858 205140 2864
rect 204168 1352 204220 1358
rect 204168 1294 204220 1300
rect 205100 480 205128 2858
rect 206204 480 206232 3062
rect 206940 3058 207506 3074
rect 206928 3052 207506 3058
rect 206980 3046 207506 3052
rect 208412 3046 208610 3074
rect 209424 3046 209714 3074
rect 206928 2994 206980 3000
rect 208412 2854 208440 3046
rect 209424 2990 209452 3046
rect 209412 2984 209464 2990
rect 209412 2926 209464 2932
rect 208400 2848 208452 2854
rect 208400 2790 208452 2796
rect 208584 2848 208636 2854
rect 208584 2790 208636 2796
rect 207388 1352 207440 1358
rect 207388 1294 207440 1300
rect 207400 480 207428 1294
rect 208596 480 208624 2790
rect 209884 1578 209912 3130
rect 211620 3120 211672 3126
rect 210528 3046 210818 3074
rect 211672 3068 211922 3074
rect 211620 3062 211922 3068
rect 210976 3052 211028 3058
rect 210528 2922 210556 3046
rect 211632 3046 211922 3062
rect 210976 2994 211028 3000
rect 210516 2916 210568 2922
rect 210516 2858 210568 2864
rect 209792 1550 209912 1578
rect 209792 480 209820 1550
rect 210988 480 211016 2994
rect 212172 2984 212224 2990
rect 212172 2926 212224 2932
rect 212184 480 212212 2926
rect 213012 1358 213040 3060
rect 213840 3046 214130 3074
rect 213368 2916 213420 2922
rect 213368 2858 213420 2864
rect 213000 1352 213052 1358
rect 213000 1294 213052 1300
rect 213380 480 213408 2858
rect 213840 2854 213868 3046
rect 213828 2848 213880 2854
rect 213828 2790 213880 2796
rect 214484 480 214512 3198
rect 214944 3194 215234 3210
rect 530032 3256 530084 3262
rect 219348 3198 219400 3204
rect 214932 3188 215234 3194
rect 214984 3182 215234 3188
rect 214932 3130 214984 3136
rect 216864 3120 216916 3126
rect 216048 3058 216338 3074
rect 219360 3074 219388 3198
rect 224880 3194 225170 3210
rect 220452 3188 220504 3194
rect 220452 3130 220504 3136
rect 224868 3188 225170 3194
rect 224920 3182 225170 3188
rect 529966 3204 530032 3210
rect 529966 3198 530084 3204
rect 546684 3256 546736 3262
rect 556712 3256 556764 3262
rect 546684 3198 546736 3204
rect 556462 3204 556712 3210
rect 556462 3198 556764 3204
rect 529966 3182 530072 3198
rect 224868 3130 224920 3136
rect 216864 3062 216916 3068
rect 216036 3052 216338 3058
rect 216088 3046 216338 3052
rect 216036 2994 216088 3000
rect 215668 2848 215720 2854
rect 215668 2790 215720 2796
rect 215680 480 215708 2790
rect 216876 480 216904 3062
rect 217152 3046 217442 3074
rect 218060 3052 218112 3058
rect 217152 2990 217180 3046
rect 218060 2994 218112 3000
rect 218256 3046 218546 3074
rect 219360 3046 219650 3074
rect 217140 2984 217192 2990
rect 217140 2926 217192 2932
rect 218072 480 218100 2994
rect 218256 2922 218284 3046
rect 218244 2916 218296 2922
rect 218244 2858 218296 2864
rect 219256 2916 219308 2922
rect 219256 2858 219308 2864
rect 219268 480 219296 2858
rect 220464 480 220492 3130
rect 221556 3120 221608 3126
rect 231032 3120 231084 3126
rect 221608 3068 221858 3074
rect 221556 3062 221858 3068
rect 220740 2854 220768 3060
rect 221568 3046 221858 3062
rect 222672 3058 222962 3074
rect 222660 3052 222962 3058
rect 222712 3046 222962 3052
rect 223500 3046 224066 3074
rect 225512 3052 225564 3058
rect 222660 2994 222712 3000
rect 222752 2984 222804 2990
rect 222752 2926 222804 2932
rect 220728 2848 220780 2854
rect 220728 2790 220780 2796
rect 221556 2848 221608 2854
rect 221556 2790 221608 2796
rect 221568 480 221596 2790
rect 222764 480 222792 2926
rect 223500 2922 223528 3046
rect 225512 2994 225564 3000
rect 223488 2916 223540 2922
rect 223488 2858 223540 2864
rect 223948 2916 224000 2922
rect 223948 2858 224000 2864
rect 223960 480 223988 2858
rect 197882 326 198320 354
rect 197882 -960 197994 326
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 354 225226 480
rect 225524 354 225552 2994
rect 226260 2854 226288 3060
rect 227364 2990 227392 3060
rect 227352 2984 227404 2990
rect 227352 2926 227404 2932
rect 227536 2984 227588 2990
rect 227536 2926 227588 2932
rect 226248 2848 226300 2854
rect 226248 2790 226300 2796
rect 226340 2848 226392 2854
rect 226340 2790 226392 2796
rect 226352 480 226380 2790
rect 227548 480 227576 2926
rect 228468 2922 228496 3060
rect 229296 3058 229586 3074
rect 234804 3120 234856 3126
rect 231032 3062 231084 3068
rect 229284 3052 229586 3058
rect 229336 3046 229586 3052
rect 229836 3052 229888 3058
rect 229284 2994 229336 3000
rect 229836 2994 229888 3000
rect 228456 2916 228508 2922
rect 228456 2858 228508 2864
rect 228732 2916 228784 2922
rect 228732 2858 228784 2864
rect 228744 480 228772 2858
rect 229848 480 229876 2994
rect 230676 2854 230704 3060
rect 230664 2848 230716 2854
rect 230664 2790 230716 2796
rect 231044 480 231072 3062
rect 231780 2990 231808 3060
rect 231768 2984 231820 2990
rect 231768 2926 231820 2932
rect 232228 2984 232280 2990
rect 232228 2926 232280 2932
rect 232240 480 232268 2926
rect 232884 2922 232912 3060
rect 233712 3058 234002 3074
rect 239312 3120 239364 3126
rect 234856 3068 235106 3074
rect 234804 3062 235106 3068
rect 233700 3052 234002 3058
rect 233752 3046 234002 3052
rect 234620 3052 234672 3058
rect 233700 2994 233752 3000
rect 234816 3046 235106 3062
rect 234620 2994 234672 3000
rect 232872 2916 232924 2922
rect 232872 2858 232924 2864
rect 233424 2848 233476 2854
rect 233424 2790 233476 2796
rect 233436 480 233464 2790
rect 234632 480 234660 2994
rect 236196 2990 236224 3060
rect 236184 2984 236236 2990
rect 236184 2926 236236 2932
rect 237012 2984 237064 2990
rect 237012 2926 237064 2932
rect 235816 2916 235868 2922
rect 235816 2858 235868 2864
rect 235828 480 235856 2858
rect 237024 480 237052 2926
rect 237300 2854 237328 3060
rect 238128 3058 238418 3074
rect 239312 3062 239364 3068
rect 242532 3120 242584 3126
rect 532608 3120 532660 3126
rect 242584 3068 242834 3074
rect 242532 3062 242834 3068
rect 238116 3052 238418 3058
rect 238168 3046 238418 3052
rect 238116 2994 238168 3000
rect 237288 2848 237340 2854
rect 237288 2790 237340 2796
rect 238116 2848 238168 2854
rect 238116 2790 238168 2796
rect 238128 480 238156 2790
rect 239324 480 239352 3062
rect 239508 2922 239536 3060
rect 240508 3052 240560 3058
rect 240508 2994 240560 3000
rect 239496 2916 239548 2922
rect 239496 2858 239548 2864
rect 240520 480 240548 2994
rect 240612 2990 240640 3060
rect 240600 2984 240652 2990
rect 240600 2926 240652 2932
rect 241716 2854 241744 3060
rect 242544 3046 242834 3062
rect 243648 3058 243938 3074
rect 243636 3052 243938 3058
rect 243688 3046 243938 3052
rect 243636 2994 243688 3000
rect 242900 2984 242952 2990
rect 242900 2926 242952 2932
rect 242072 2916 242124 2922
rect 242072 2858 242124 2864
rect 241704 2848 241756 2854
rect 241704 2790 241756 2796
rect 225114 326 225552 354
rect 225114 -960 225226 326
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 354 241786 480
rect 242084 354 242112 2858
rect 242912 480 242940 2926
rect 245028 2922 245056 3060
rect 246132 2990 246160 3060
rect 246120 2984 246172 2990
rect 246120 2926 246172 2932
rect 246396 2984 246448 2990
rect 246396 2926 246448 2932
rect 245016 2916 245068 2922
rect 245016 2858 245068 2864
rect 245200 2916 245252 2922
rect 245200 2858 245252 2864
rect 244096 2848 244148 2854
rect 244096 2790 244148 2796
rect 244108 480 244136 2790
rect 245212 480 245240 2858
rect 246408 480 246436 2926
rect 247236 2854 247264 3060
rect 248340 2922 248368 3060
rect 248788 3052 248840 3058
rect 248788 2994 248840 3000
rect 248328 2916 248380 2922
rect 248328 2858 248380 2864
rect 247224 2848 247276 2854
rect 247224 2790 247276 2796
rect 247592 2848 247644 2854
rect 247592 2790 247644 2796
rect 247604 480 247632 2790
rect 248800 480 248828 2994
rect 249444 2990 249472 3060
rect 249432 2984 249484 2990
rect 249432 2926 249484 2932
rect 249984 2916 250036 2922
rect 249984 2858 250036 2864
rect 249996 480 250024 2858
rect 250548 2854 250576 3060
rect 251376 3058 251666 3074
rect 251364 3052 251666 3058
rect 251416 3046 251666 3052
rect 251364 2994 251416 3000
rect 252756 2922 252784 3060
rect 253480 2984 253532 2990
rect 253480 2926 253532 2932
rect 252744 2916 252796 2922
rect 252744 2858 252796 2864
rect 250536 2848 250588 2854
rect 250536 2790 250588 2796
rect 252376 2848 252428 2854
rect 252376 2790 252428 2796
rect 251180 808 251232 814
rect 251180 750 251232 756
rect 251192 480 251220 750
rect 252388 480 252416 2790
rect 253492 480 253520 2926
rect 253860 814 253888 3060
rect 254676 2916 254728 2922
rect 254676 2858 254728 2864
rect 253848 808 253900 814
rect 253848 750 253900 756
rect 254688 480 254716 2858
rect 254964 2854 254992 3060
rect 256068 2990 256096 3060
rect 256056 2984 256108 2990
rect 256056 2926 256108 2932
rect 257172 2922 257200 3060
rect 257160 2916 257212 2922
rect 257160 2858 257212 2864
rect 258276 2854 258304 3060
rect 254952 2848 255004 2854
rect 254952 2790 255004 2796
rect 255872 2848 255924 2854
rect 255872 2790 255924 2796
rect 258264 2848 258316 2854
rect 258264 2790 258316 2796
rect 255884 480 255912 2790
rect 259380 1358 259408 3060
rect 257068 1352 257120 1358
rect 257068 1294 257120 1300
rect 259368 1352 259420 1358
rect 259368 1294 259420 1300
rect 259460 1352 259512 1358
rect 259460 1294 259512 1300
rect 257080 480 257108 1294
rect 258264 1284 258316 1290
rect 258264 1226 258316 1232
rect 258276 480 258304 1226
rect 259472 480 259500 1294
rect 260484 1290 260512 3060
rect 260656 2848 260708 2854
rect 260656 2790 260708 2796
rect 260472 1284 260524 1290
rect 260472 1226 260524 1232
rect 260668 480 260696 2790
rect 261588 1358 261616 3060
rect 261760 2916 261812 2922
rect 261760 2858 261812 2864
rect 261576 1352 261628 1358
rect 261576 1294 261628 1300
rect 261772 480 261800 2858
rect 262692 2854 262720 3060
rect 263796 2922 263824 3060
rect 263784 2916 263836 2922
rect 263784 2858 263836 2864
rect 262680 2848 262732 2854
rect 262680 2790 262732 2796
rect 264900 1358 264928 3060
rect 262956 1352 263008 1358
rect 262956 1294 263008 1300
rect 264888 1352 264940 1358
rect 264888 1294 264940 1300
rect 265348 1352 265400 1358
rect 265348 1294 265400 1300
rect 262968 480 262996 1294
rect 264152 1284 264204 1290
rect 264152 1226 264204 1232
rect 264164 480 264192 1226
rect 265360 480 265388 1294
rect 266004 1290 266032 3060
rect 267108 1358 267136 3060
rect 267096 1352 267148 1358
rect 267096 1294 267148 1300
rect 267740 1352 267792 1358
rect 267740 1294 267792 1300
rect 265992 1284 266044 1290
rect 265992 1226 266044 1232
rect 266544 1284 266596 1290
rect 266544 1226 266596 1232
rect 266556 480 266584 1226
rect 267752 480 267780 1294
rect 268212 1290 268240 3060
rect 269316 1358 269344 3060
rect 269304 1352 269356 1358
rect 269304 1294 269356 1300
rect 268200 1284 268252 1290
rect 268200 1226 268252 1232
rect 270040 1284 270092 1290
rect 270040 1226 270092 1232
rect 268844 1216 268896 1222
rect 268844 1158 268896 1164
rect 268856 480 268884 1158
rect 270052 480 270080 1226
rect 270420 1222 270448 3060
rect 271236 1352 271288 1358
rect 271236 1294 271288 1300
rect 270408 1216 270460 1222
rect 270408 1158 270460 1164
rect 271248 480 271276 1294
rect 271524 1290 271552 3060
rect 272628 1358 272656 3060
rect 272616 1352 272668 1358
rect 272616 1294 272668 1300
rect 273628 1352 273680 1358
rect 273628 1294 273680 1300
rect 271512 1284 271564 1290
rect 271512 1226 271564 1232
rect 272432 1284 272484 1290
rect 272432 1226 272484 1232
rect 272444 480 272472 1226
rect 273640 480 273668 1294
rect 273732 1290 273760 3060
rect 274836 1358 274864 3060
rect 275296 3046 275954 3074
rect 276124 3046 277058 3074
rect 274824 1352 274876 1358
rect 274824 1294 274876 1300
rect 273720 1284 273772 1290
rect 273720 1226 273772 1232
rect 241674 326 242112 354
rect 241674 -960 241786 326
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 354 274906 480
rect 275296 354 275324 3046
rect 276124 1578 276152 3046
rect 276032 1550 276152 1578
rect 276032 480 276060 1550
rect 278148 1358 278176 3060
rect 278792 3046 279266 3074
rect 277124 1352 277176 1358
rect 277124 1294 277176 1300
rect 278136 1352 278188 1358
rect 278136 1294 278188 1300
rect 277136 480 277164 1294
rect 274794 326 275324 354
rect 274794 -960 274906 326
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 354 278402 480
rect 278792 354 278820 3046
rect 280356 1358 280384 3060
rect 281184 3046 281474 3074
rect 281920 3046 282578 3074
rect 283392 3046 283682 3074
rect 284312 3046 284786 3074
rect 285416 3046 285890 3074
rect 279516 1352 279568 1358
rect 279516 1294 279568 1300
rect 280344 1352 280396 1358
rect 280344 1294 280396 1300
rect 279528 480 279556 1294
rect 278290 326 278820 354
rect 278290 -960 278402 326
rect 279486 -960 279598 480
rect 280682 354 280794 480
rect 281184 354 281212 3046
rect 281920 480 281948 3046
rect 280682 326 281212 354
rect 280682 -960 280794 326
rect 281878 -960 281990 480
rect 283074 354 283186 480
rect 283392 354 283420 3046
rect 284312 480 284340 3046
rect 285416 480 285444 3046
rect 283074 326 283420 354
rect 283074 -960 283186 326
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 354 286682 480
rect 286980 354 287008 3060
rect 287808 3046 288098 3074
rect 287808 480 287836 3046
rect 286570 326 287008 354
rect 286570 -960 286682 326
rect 287766 -960 287878 480
rect 288962 354 289074 480
rect 289188 354 289216 3060
rect 290200 3046 290306 3074
rect 290200 480 290228 3046
rect 291396 480 291424 3060
rect 292592 480 292620 3060
rect 293696 480 293724 3060
rect 294814 3046 294920 3074
rect 295918 3046 296116 3074
rect 297022 3046 297312 3074
rect 294892 480 294920 3046
rect 296088 480 296116 3046
rect 297284 480 297312 3046
rect 288962 326 289216 354
rect 288962 -960 289074 326
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298112 354 298140 3060
rect 299230 3046 299704 3074
rect 300334 3046 300808 3074
rect 301438 3046 301728 3074
rect 302542 3046 303200 3074
rect 303646 3046 303936 3074
rect 299676 480 299704 3046
rect 300780 480 300808 3046
rect 298438 354 298550 480
rect 298112 326 298550 354
rect 298438 -960 298550 326
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301700 354 301728 3046
rect 303172 480 303200 3046
rect 301934 354 302046 480
rect 301700 326 302046 354
rect 301934 -960 302046 326
rect 303130 -960 303242 480
rect 303908 354 303936 3046
rect 304736 2854 304764 3060
rect 305854 3046 306328 3074
rect 304724 2848 304776 2854
rect 304724 2790 304776 2796
rect 305552 2848 305604 2854
rect 305552 2790 305604 2796
rect 305564 480 305592 2790
rect 304326 354 304438 480
rect 303908 326 304438 354
rect 304326 -960 304438 326
rect 305522 -960 305634 480
rect 306300 354 306328 3046
rect 306944 2854 306972 3060
rect 308062 3046 308996 3074
rect 306932 2848 306984 2854
rect 306932 2790 306984 2796
rect 307944 2848 307996 2854
rect 307944 2790 307996 2796
rect 307956 480 307984 2790
rect 308968 1578 308996 3046
rect 309152 2854 309180 3060
rect 310256 2990 310284 3060
rect 310244 2984 310296 2990
rect 310244 2926 310296 2932
rect 311360 2854 311388 3060
rect 311440 2984 311492 2990
rect 311440 2926 311492 2932
rect 309140 2848 309192 2854
rect 309140 2790 309192 2796
rect 310244 2848 310296 2854
rect 310244 2790 310296 2796
rect 311348 2848 311400 2854
rect 311348 2790 311400 2796
rect 308968 1550 309088 1578
rect 309060 480 309088 1550
rect 310256 480 310284 2790
rect 311452 480 311480 2926
rect 312464 2922 312492 3060
rect 312452 2916 312504 2922
rect 312452 2858 312504 2864
rect 313568 2854 313596 3060
rect 314580 2922 314608 3060
rect 313832 2916 313884 2922
rect 313832 2858 313884 2864
rect 314568 2916 314620 2922
rect 314568 2858 314620 2864
rect 312636 2848 312688 2854
rect 312636 2790 312688 2796
rect 313556 2848 313608 2854
rect 313556 2790 313608 2796
rect 312648 480 312676 2790
rect 313844 480 313872 2858
rect 315776 2854 315804 3060
rect 316880 2922 316908 3060
rect 316224 2916 316276 2922
rect 316224 2858 316276 2864
rect 316868 2916 316920 2922
rect 316868 2858 316920 2864
rect 315028 2848 315080 2854
rect 315028 2790 315080 2796
rect 315764 2848 315816 2854
rect 315764 2790 315816 2796
rect 315040 480 315068 2790
rect 316236 480 316264 2858
rect 317984 2854 318012 3060
rect 319088 2922 319116 3060
rect 318524 2916 318576 2922
rect 318524 2858 318576 2864
rect 319076 2916 319128 2922
rect 319076 2858 319128 2864
rect 317328 2848 317380 2854
rect 317328 2790 317380 2796
rect 317972 2848 318024 2854
rect 317972 2790 318024 2796
rect 317340 480 317368 2790
rect 318536 480 318564 2858
rect 320100 2854 320128 3060
rect 321296 2922 321324 3060
rect 320916 2916 320968 2922
rect 320916 2858 320968 2864
rect 321284 2916 321336 2922
rect 321284 2858 321336 2864
rect 319720 2848 319772 2854
rect 319720 2790 319772 2796
rect 320088 2848 320140 2854
rect 320088 2790 320140 2796
rect 319732 480 319760 2790
rect 320928 480 320956 2858
rect 322400 2854 322428 3060
rect 323504 2922 323532 3060
rect 323308 2916 323360 2922
rect 323308 2858 323360 2864
rect 323492 2916 323544 2922
rect 323492 2858 323544 2864
rect 322112 2848 322164 2854
rect 322112 2790 322164 2796
rect 322388 2848 322440 2854
rect 322388 2790 322440 2796
rect 322124 480 322152 2790
rect 323320 480 323348 2858
rect 324608 2854 324636 3060
rect 325712 2990 325740 3060
rect 326830 3046 327028 3074
rect 325700 2984 325752 2990
rect 325700 2926 325752 2932
rect 325608 2916 325660 2922
rect 325608 2858 325660 2864
rect 324412 2848 324464 2854
rect 324412 2790 324464 2796
rect 324596 2848 324648 2854
rect 324596 2790 324648 2796
rect 324424 480 324452 2790
rect 325620 480 325648 2858
rect 327000 2854 327028 3046
rect 327920 2922 327948 3060
rect 329024 2990 329052 3060
rect 328000 2984 328052 2990
rect 328000 2926 328052 2932
rect 329012 2984 329064 2990
rect 329012 2926 329064 2932
rect 327908 2916 327960 2922
rect 327908 2858 327960 2864
rect 326804 2848 326856 2854
rect 326804 2790 326856 2796
rect 326988 2848 327040 2854
rect 326988 2790 327040 2796
rect 326816 480 326844 2790
rect 328012 480 328040 2926
rect 330128 2854 330156 3060
rect 331246 3058 331352 3074
rect 331246 3052 331364 3058
rect 331246 3046 331312 3052
rect 331312 2994 331364 3000
rect 332336 2990 332364 3060
rect 331588 2984 331640 2990
rect 331588 2926 331640 2932
rect 332324 2984 332376 2990
rect 332324 2926 332376 2932
rect 330392 2916 330444 2922
rect 330392 2858 330444 2864
rect 329196 2848 329248 2854
rect 329196 2790 329248 2796
rect 330116 2848 330168 2854
rect 330116 2790 330168 2796
rect 329208 480 329236 2790
rect 330404 480 330432 2858
rect 331600 480 331628 2926
rect 333440 2922 333468 3060
rect 334558 3058 334848 3074
rect 333888 3052 333940 3058
rect 334558 3052 334860 3058
rect 334558 3046 334808 3052
rect 333888 2994 333940 3000
rect 334808 2994 334860 3000
rect 333428 2916 333480 2922
rect 333428 2858 333480 2864
rect 332692 2848 332744 2854
rect 332692 2790 332744 2796
rect 332704 480 332732 2790
rect 333900 480 333928 2994
rect 335084 2984 335136 2990
rect 335084 2926 335136 2932
rect 335096 480 335124 2926
rect 335648 2854 335676 3060
rect 336280 2916 336332 2922
rect 336280 2858 336332 2864
rect 335636 2848 335688 2854
rect 335636 2790 335688 2796
rect 336292 480 336320 2858
rect 336660 1358 336688 3060
rect 337476 3052 337528 3058
rect 337476 2994 337528 3000
rect 336648 1352 336700 1358
rect 336648 1294 336700 1300
rect 337488 480 337516 2994
rect 337856 882 337884 3060
rect 338960 2854 338988 3060
rect 340064 2922 340092 3060
rect 341168 2990 341196 3060
rect 341156 2984 341208 2990
rect 341156 2926 341208 2932
rect 340052 2916 340104 2922
rect 340052 2858 340104 2864
rect 338672 2848 338724 2854
rect 338672 2790 338724 2796
rect 338948 2848 339000 2854
rect 338948 2790 339000 2796
rect 342076 2848 342128 2854
rect 342076 2790 342128 2796
rect 337844 876 337896 882
rect 337844 818 337896 824
rect 338684 480 338712 2790
rect 339868 1352 339920 1358
rect 339868 1294 339920 1300
rect 339880 480 339908 1294
rect 342088 1170 342116 2790
rect 342180 1358 342208 3060
rect 342996 2916 343048 2922
rect 342996 2858 343048 2864
rect 342168 1352 342220 1358
rect 342168 1294 342220 1300
rect 342088 1142 342208 1170
rect 340972 876 341024 882
rect 340972 818 341024 824
rect 340984 480 341012 818
rect 342180 480 342208 1142
rect 306718 354 306830 480
rect 306300 326 306830 354
rect 306718 -960 306830 326
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343008 354 343036 2858
rect 343376 1290 343404 3060
rect 344494 3046 344784 3074
rect 344560 2984 344612 2990
rect 344560 2926 344612 2932
rect 343364 1284 343416 1290
rect 343364 1226 343416 1232
rect 344572 480 344600 2926
rect 343334 354 343446 480
rect 343008 326 343446 354
rect 343334 -960 343446 326
rect 344530 -960 344642 480
rect 344756 66 344784 3046
rect 345584 1018 345612 3060
rect 346688 2854 346716 3060
rect 346676 2848 346728 2854
rect 346676 2790 346728 2796
rect 345756 1352 345808 1358
rect 345756 1294 345808 1300
rect 345572 1012 345624 1018
rect 345572 954 345624 960
rect 345768 480 345796 1294
rect 346952 1284 347004 1290
rect 346952 1226 347004 1232
rect 346964 480 346992 1226
rect 347700 882 347728 3060
rect 348896 1358 348924 3060
rect 348884 1352 348936 1358
rect 348884 1294 348936 1300
rect 350000 1290 350028 3060
rect 350448 2848 350500 2854
rect 350448 2790 350500 2796
rect 349988 1284 350040 1290
rect 349988 1226 350040 1232
rect 349252 1012 349304 1018
rect 349252 954 349304 960
rect 347688 876 347740 882
rect 347688 818 347740 824
rect 349264 480 349292 954
rect 350460 480 350488 2790
rect 351104 1018 351132 3060
rect 352208 1154 352236 3060
rect 353220 2854 353248 3060
rect 353208 2848 353260 2854
rect 353208 2790 353260 2796
rect 352840 1352 352892 1358
rect 352840 1294 352892 1300
rect 352196 1148 352248 1154
rect 352196 1090 352248 1096
rect 351092 1012 351144 1018
rect 351092 954 351144 960
rect 351644 876 351696 882
rect 351644 818 351696 824
rect 351656 480 351684 818
rect 352852 480 352880 1294
rect 354036 1284 354088 1290
rect 354036 1226 354088 1232
rect 354048 480 354076 1226
rect 344744 60 344796 66
rect 344744 2 344796 8
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 82 348138 480
rect 348026 66 348280 82
rect 348026 60 348292 66
rect 348026 54 348240 60
rect 348026 -960 348138 54
rect 348240 2 348292 8
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 354416 134 354444 3060
rect 355520 1086 355548 3060
rect 356624 1358 356652 3060
rect 357532 2848 357584 2854
rect 357532 2790 357584 2796
rect 356612 1352 356664 1358
rect 356612 1294 356664 1300
rect 356336 1148 356388 1154
rect 356336 1090 356388 1096
rect 355508 1080 355560 1086
rect 355508 1022 355560 1028
rect 355232 1012 355284 1018
rect 355232 954 355284 960
rect 355244 480 355272 954
rect 356348 480 356376 1090
rect 357544 480 357572 2790
rect 357728 1290 357756 3060
rect 357716 1284 357768 1290
rect 357716 1226 357768 1232
rect 358740 950 358768 3060
rect 359936 1222 359964 3060
rect 359924 1216 359976 1222
rect 359924 1158 359976 1164
rect 361040 1154 361068 3060
rect 361120 1352 361172 1358
rect 361120 1294 361172 1300
rect 361028 1148 361080 1154
rect 361028 1090 361080 1096
rect 359924 1080 359976 1086
rect 359924 1022 359976 1028
rect 358728 944 358780 950
rect 358728 886 358780 892
rect 359936 480 359964 1022
rect 361132 480 361160 1294
rect 362144 1018 362172 3060
rect 362316 1284 362368 1290
rect 362316 1226 362368 1232
rect 362132 1012 362184 1018
rect 362132 954 362184 960
rect 362328 480 362356 1226
rect 354404 128 354456 134
rect 354404 70 354456 76
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 82 358810 480
rect 358912 128 358964 134
rect 358698 76 358912 82
rect 358698 70 358964 76
rect 358698 54 358952 70
rect 358698 -960 358810 54
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363248 134 363276 3060
rect 364260 1358 364288 3060
rect 364248 1352 364300 1358
rect 364248 1294 364300 1300
rect 365456 1290 365484 3060
rect 365444 1284 365496 1290
rect 365444 1226 365496 1232
rect 364616 1216 364668 1222
rect 364616 1158 364668 1164
rect 363512 944 363564 950
rect 363512 886 363564 892
rect 363524 480 363552 886
rect 364628 480 364656 1158
rect 365444 1148 365496 1154
rect 365444 1090 365496 1096
rect 363236 128 363288 134
rect 363236 70 363288 76
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365456 354 365484 1090
rect 366560 1086 366588 3060
rect 366548 1080 366600 1086
rect 366548 1022 366600 1028
rect 367664 1018 367692 3060
rect 368768 1222 368796 3060
rect 369400 1352 369452 1358
rect 369400 1294 369452 1300
rect 368756 1216 368808 1222
rect 368756 1158 368808 1164
rect 367008 1012 367060 1018
rect 367008 954 367060 960
rect 367652 1012 367704 1018
rect 367652 954 367704 960
rect 367020 480 367048 954
rect 369412 480 369440 1294
rect 369780 1154 369808 3060
rect 370976 1290 371004 3060
rect 372094 3046 372384 3074
rect 372356 2854 372384 3046
rect 372344 2848 372396 2854
rect 372344 2790 372396 2796
rect 370228 1284 370280 1290
rect 370228 1226 370280 1232
rect 370964 1284 371016 1290
rect 370964 1226 371016 1232
rect 369768 1148 369820 1154
rect 369768 1090 369820 1096
rect 365782 354 365894 480
rect 365456 326 365894 354
rect 365782 -960 365894 326
rect 366978 -960 367090 480
rect 367836 128 367888 134
rect 368174 82 368286 480
rect 367888 76 368286 82
rect 367836 70 368286 76
rect 367848 54 368286 70
rect 368174 -960 368286 54
rect 369370 -960 369482 480
rect 370240 354 370268 1226
rect 373184 1086 373212 3060
rect 374288 1358 374316 3060
rect 375208 3046 375314 3074
rect 374276 1352 374328 1358
rect 374276 1294 374328 1300
rect 373908 1216 373960 1222
rect 373908 1158 373960 1164
rect 371332 1080 371384 1086
rect 371332 1022 371384 1028
rect 373172 1080 373224 1086
rect 373172 1022 373224 1028
rect 370566 354 370678 480
rect 370240 326 370678 354
rect 371344 354 371372 1022
rect 372896 1012 372948 1018
rect 372896 954 372948 960
rect 372908 480 372936 954
rect 371670 354 371782 480
rect 371344 326 371782 354
rect 370566 -960 370678 326
rect 371670 -960 371782 326
rect 372866 -960 372978 480
rect 373920 354 373948 1158
rect 375208 1018 375236 3046
rect 376496 1290 376524 3060
rect 376116 1284 376168 1290
rect 376116 1226 376168 1232
rect 376484 1284 376536 1290
rect 376484 1226 376536 1232
rect 375288 1148 375340 1154
rect 375288 1090 375340 1096
rect 375196 1012 375248 1018
rect 375196 954 375248 960
rect 375300 480 375328 1090
rect 374062 354 374174 480
rect 373920 326 374174 354
rect 374062 -960 374174 326
rect 375258 -960 375370 480
rect 376128 354 376156 1226
rect 377600 950 377628 3060
rect 377680 2848 377732 2854
rect 377680 2790 377732 2796
rect 377588 944 377640 950
rect 377588 886 377640 892
rect 377692 480 377720 2790
rect 378704 1222 378732 3060
rect 379612 1352 379664 1358
rect 379612 1294 379664 1300
rect 378692 1216 378744 1222
rect 378692 1158 378744 1164
rect 378508 1080 378560 1086
rect 378508 1022 378560 1028
rect 376454 354 376566 480
rect 376128 326 376566 354
rect 376454 -960 376566 326
rect 377650 -960 377762 480
rect 378520 354 378548 1022
rect 378846 354 378958 480
rect 378520 326 378958 354
rect 379624 354 379652 1294
rect 379808 1154 379836 3060
rect 379796 1148 379848 1154
rect 379796 1090 379848 1096
rect 379950 354 380062 480
rect 379624 326 380062 354
rect 378846 -960 378958 326
rect 379950 -960 380062 326
rect 380820 270 380848 3060
rect 381176 1012 381228 1018
rect 381176 954 381228 960
rect 381188 480 381216 954
rect 380808 264 380860 270
rect 380808 206 380860 212
rect 381146 -960 381258 480
rect 382016 474 382044 3060
rect 382372 1284 382424 1290
rect 382372 1226 382424 1232
rect 382384 480 382412 1226
rect 382004 468 382056 474
rect 382004 410 382056 416
rect 382342 -960 382454 480
rect 383120 66 383148 3060
rect 383568 944 383620 950
rect 383568 886 383620 892
rect 383580 480 383608 886
rect 384224 610 384252 3060
rect 385328 1358 385356 3060
rect 385316 1352 385368 1358
rect 385316 1294 385368 1300
rect 384396 1216 384448 1222
rect 384396 1158 384448 1164
rect 384212 604 384264 610
rect 384212 546 384264 552
rect 383108 60 383160 66
rect 383108 2 383160 8
rect 383538 -960 383650 480
rect 384408 354 384436 1158
rect 385960 1148 386012 1154
rect 385960 1090 386012 1096
rect 385972 480 386000 1090
rect 386340 882 386368 3060
rect 387536 1222 387564 3060
rect 388640 1290 388668 3060
rect 388628 1284 388680 1290
rect 388628 1226 388680 1232
rect 387524 1216 387576 1222
rect 387524 1158 387576 1164
rect 386328 876 386380 882
rect 386328 818 386380 824
rect 384734 354 384846 480
rect 384408 326 384846 354
rect 384734 -960 384846 326
rect 385930 -960 386042 480
rect 386788 264 386840 270
rect 387126 218 387238 480
rect 387892 468 387944 474
rect 387892 410 387944 416
rect 387904 354 387932 410
rect 388230 354 388342 480
rect 387904 326 388342 354
rect 386840 212 387238 218
rect 386788 206 387238 212
rect 386800 190 387238 206
rect 387126 -960 387238 190
rect 388230 -960 388342 326
rect 389426 82 389538 480
rect 389744 202 389772 3060
rect 390652 604 390704 610
rect 390652 546 390704 552
rect 390664 480 390692 546
rect 390848 542 390876 3060
rect 391676 3046 391874 3074
rect 390836 536 390888 542
rect 389732 196 389784 202
rect 389732 138 389784 144
rect 389426 66 389680 82
rect 389426 60 389692 66
rect 389426 54 389640 60
rect 389426 -960 389538 54
rect 389640 2 389692 8
rect 390622 -960 390734 480
rect 390836 478 390888 484
rect 391676 338 391704 3046
rect 391848 1352 391900 1358
rect 391848 1294 391900 1300
rect 391860 480 391888 1294
rect 392676 876 392728 882
rect 392676 818 392728 824
rect 391664 332 391716 338
rect 391664 274 391716 280
rect 391818 -960 391930 480
rect 392688 218 392716 818
rect 393056 610 393084 3060
rect 394160 1086 394188 3060
rect 395264 1222 395292 3060
rect 396368 1358 396396 3060
rect 396356 1352 396408 1358
rect 396356 1294 396408 1300
rect 395344 1284 395396 1290
rect 395344 1226 395396 1232
rect 394240 1216 394292 1222
rect 394240 1158 394292 1164
rect 395252 1216 395304 1222
rect 395252 1158 395304 1164
rect 394148 1080 394200 1086
rect 394148 1022 394200 1028
rect 393044 604 393096 610
rect 393044 546 393096 552
rect 394252 480 394280 1158
rect 395356 480 395384 1226
rect 397380 1154 397408 3060
rect 397368 1148 397420 1154
rect 397368 1090 397420 1096
rect 397736 604 397788 610
rect 397736 546 397788 552
rect 397748 480 397776 546
rect 393014 218 393126 480
rect 392688 190 393126 218
rect 393014 -960 393126 190
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 218 396622 480
rect 396184 202 396622 218
rect 396172 196 396622 202
rect 396224 190 396622 196
rect 396172 138 396224 144
rect 396510 -960 396622 190
rect 397706 -960 397818 480
rect 398576 270 398604 3060
rect 398902 354 399014 480
rect 398760 338 399014 354
rect 398748 332 399014 338
rect 398800 326 399014 332
rect 398748 274 398800 280
rect 398564 264 398616 270
rect 398564 206 398616 212
rect 398902 -960 399014 326
rect 399680 202 399708 3060
rect 400128 672 400180 678
rect 400128 614 400180 620
rect 400140 480 400168 614
rect 399668 196 399720 202
rect 399668 138 399720 144
rect 400098 -960 400210 480
rect 400784 338 400812 3060
rect 401324 1080 401376 1086
rect 401324 1022 401376 1028
rect 401336 480 401364 1022
rect 401888 678 401916 3060
rect 402520 1216 402572 1222
rect 402520 1158 402572 1164
rect 401876 672 401928 678
rect 401876 614 401928 620
rect 402532 480 402560 1158
rect 400772 332 400824 338
rect 400772 274 400824 280
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 402900 134 402928 3060
rect 403624 1352 403676 1358
rect 403624 1294 403676 1300
rect 403636 480 403664 1294
rect 404096 1290 404124 3060
rect 404084 1284 404136 1290
rect 404084 1226 404136 1232
rect 404820 1148 404872 1154
rect 404820 1090 404872 1096
rect 404832 480 404860 1090
rect 402888 128 402940 134
rect 402888 70 402940 76
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405200 406 405228 3060
rect 406304 1358 406332 3060
rect 406292 1352 406344 1358
rect 406292 1294 406344 1300
rect 405188 400 405240 406
rect 405188 342 405240 348
rect 405986 218 406098 480
rect 406200 264 406252 270
rect 405986 212 406200 218
rect 407182 218 407294 480
rect 405986 206 406252 212
rect 405986 190 406240 206
rect 407040 202 407294 218
rect 407408 202 407436 3060
rect 408420 610 408448 3060
rect 409236 672 409288 678
rect 409236 614 409288 620
rect 408408 604 408460 610
rect 408408 546 408460 552
rect 408378 354 408490 480
rect 408378 338 408632 354
rect 408378 332 408644 338
rect 408378 326 408592 332
rect 407028 196 407294 202
rect 405986 -960 406098 190
rect 407080 190 407294 196
rect 407028 138 407080 144
rect 407182 -960 407294 190
rect 407396 196 407448 202
rect 407396 138 407448 144
rect 408378 -960 408490 326
rect 408592 274 408644 280
rect 409248 218 409276 614
rect 409616 610 409644 3060
rect 410734 3046 411024 3074
rect 411838 3046 412128 3074
rect 409604 604 409656 610
rect 409604 546 409656 552
rect 409574 218 409686 480
rect 409248 190 409686 218
rect 409574 -960 409686 190
rect 410770 82 410882 480
rect 410996 270 411024 3046
rect 411904 1284 411956 1290
rect 411904 1226 411956 1232
rect 411916 480 411944 1226
rect 410984 264 411036 270
rect 410984 206 411036 212
rect 410984 128 411036 134
rect 410770 76 410984 82
rect 410770 70 411036 76
rect 410770 54 411024 70
rect 410770 -960 410882 54
rect 411874 -960 411986 480
rect 412100 338 412128 3046
rect 412928 1154 412956 3060
rect 413940 1290 413968 3060
rect 415136 1358 415164 3060
rect 414296 1352 414348 1358
rect 414296 1294 414348 1300
rect 415124 1352 415176 1358
rect 415124 1294 415176 1300
rect 413928 1284 413980 1290
rect 413928 1226 413980 1232
rect 412916 1148 412968 1154
rect 412916 1090 412968 1096
rect 414308 480 414336 1294
rect 416240 950 416268 3060
rect 416228 944 416280 950
rect 416228 886 416280 892
rect 416688 604 416740 610
rect 416688 546 416740 552
rect 416700 480 416728 546
rect 412824 400 412876 406
rect 413070 354 413182 480
rect 412876 348 413182 354
rect 412824 342 413182 348
rect 412088 332 412140 338
rect 412836 326 413182 342
rect 412088 274 412140 280
rect 413070 -960 413182 326
rect 414266 -960 414378 480
rect 415462 218 415574 480
rect 415320 202 415574 218
rect 415308 196 415574 202
rect 415360 190 415574 196
rect 415308 138 415360 144
rect 415462 -960 415574 190
rect 416658 -960 416770 480
rect 417344 202 417372 3060
rect 417884 672 417936 678
rect 417884 614 417936 620
rect 417896 480 417924 614
rect 417332 196 417384 202
rect 417332 138 417384 144
rect 417854 -960 417966 480
rect 418448 406 418476 3060
rect 419460 1018 419488 3060
rect 420656 1222 420684 3060
rect 420644 1216 420696 1222
rect 420644 1158 420696 1164
rect 421380 1148 421432 1154
rect 421380 1090 421432 1096
rect 419448 1012 419500 1018
rect 419448 954 419500 960
rect 421392 480 421420 1090
rect 421760 882 421788 3060
rect 422576 1284 422628 1290
rect 422576 1226 422628 1232
rect 421748 876 421800 882
rect 421748 818 421800 824
rect 422588 480 422616 1226
rect 422864 1154 422892 3060
rect 423404 1352 423456 1358
rect 423404 1294 423456 1300
rect 422852 1148 422904 1154
rect 422852 1090 422904 1096
rect 418436 400 418488 406
rect 418436 342 418488 348
rect 418620 264 418672 270
rect 418958 218 419070 480
rect 418672 212 419070 218
rect 418620 206 419070 212
rect 418632 190 419070 206
rect 418958 -960 419070 190
rect 420154 354 420266 480
rect 420154 338 420408 354
rect 420154 332 420420 338
rect 420154 326 420368 332
rect 420154 -960 420266 326
rect 420368 274 420420 280
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423416 354 423444 1294
rect 423742 354 423854 480
rect 423416 326 423854 354
rect 423742 -960 423854 326
rect 423968 66 423996 3060
rect 424980 1086 425008 3060
rect 426176 1290 426204 3060
rect 426164 1284 426216 1290
rect 426164 1226 426216 1232
rect 424968 1080 425020 1086
rect 424968 1022 425020 1028
rect 424968 944 425020 950
rect 424968 886 425020 892
rect 424980 480 425008 886
rect 427280 678 427308 3060
rect 428384 1358 428412 3060
rect 428372 1352 428424 1358
rect 428372 1294 428424 1300
rect 429292 1216 429344 1222
rect 429292 1158 429344 1164
rect 428464 1012 428516 1018
rect 428464 954 428516 960
rect 427268 672 427320 678
rect 427268 614 427320 620
rect 428476 480 428504 954
rect 423956 60 424008 66
rect 423956 2 424008 8
rect 424938 -960 425050 480
rect 426134 218 426246 480
rect 426900 400 426952 406
rect 427238 354 427350 480
rect 426952 348 427350 354
rect 426900 342 427350 348
rect 426912 326 427350 342
rect 425808 202 426246 218
rect 425796 196 426246 202
rect 425848 190 426246 196
rect 425796 138 425848 144
rect 426134 -960 426246 190
rect 427238 -960 427350 326
rect 428434 -960 428546 480
rect 429304 354 429332 1158
rect 429488 814 429516 3060
rect 430500 950 430528 3060
rect 431696 1018 431724 3060
rect 431868 1148 431920 1154
rect 431868 1090 431920 1096
rect 431684 1012 431736 1018
rect 431684 954 431736 960
rect 430488 944 430540 950
rect 430488 886 430540 892
rect 430856 876 430908 882
rect 430856 818 430908 824
rect 429476 808 429528 814
rect 429476 750 429528 756
rect 430868 480 430896 818
rect 429630 354 429742 480
rect 429304 326 429742 354
rect 429630 -960 429742 326
rect 430826 -960 430938 480
rect 431880 354 431908 1090
rect 432800 746 432828 3060
rect 432788 740 432840 746
rect 432788 682 432840 688
rect 433904 610 433932 3060
rect 435008 1222 435036 3060
rect 436020 1290 436048 3060
rect 435180 1284 435232 1290
rect 435180 1226 435232 1232
rect 436008 1284 436060 1290
rect 436008 1226 436060 1232
rect 434996 1216 435048 1222
rect 434996 1158 435048 1164
rect 434076 1080 434128 1086
rect 434076 1022 434128 1028
rect 433892 604 433944 610
rect 433892 546 433944 552
rect 432022 354 432134 480
rect 431880 326 432134 354
rect 432022 -960 432134 326
rect 433218 82 433330 480
rect 434088 354 434116 1022
rect 434414 354 434526 480
rect 434088 326 434526 354
rect 435192 354 435220 1226
rect 437216 950 437244 3060
rect 437572 1352 437624 1358
rect 437572 1294 437624 1300
rect 437204 944 437256 950
rect 437204 886 437256 892
rect 436744 672 436796 678
rect 436744 614 436796 620
rect 436756 480 436784 614
rect 435518 354 435630 480
rect 435192 326 435630 354
rect 433218 66 433472 82
rect 433218 60 433484 66
rect 433218 54 433432 60
rect 433218 -960 433330 54
rect 433432 2 433484 8
rect 434414 -960 434526 326
rect 435518 -960 435630 326
rect 436714 -960 436826 480
rect 437584 354 437612 1294
rect 438320 1154 438348 3060
rect 439424 1358 439452 3060
rect 439412 1352 439464 1358
rect 439412 1294 439464 1300
rect 438308 1148 438360 1154
rect 438308 1090 438360 1096
rect 440332 876 440384 882
rect 440332 818 440384 824
rect 439136 808 439188 814
rect 439136 750 439188 756
rect 439148 480 439176 750
rect 440344 480 440372 818
rect 440528 814 440556 3060
rect 441540 1018 441568 3060
rect 442736 1086 442764 3060
rect 443736 1352 443788 1358
rect 443736 1294 443788 1300
rect 442724 1080 442776 1086
rect 442724 1022 442776 1028
rect 441436 1012 441488 1018
rect 441436 954 441488 960
rect 441528 1012 441580 1018
rect 441528 954 441580 960
rect 440516 808 440568 814
rect 440516 750 440568 756
rect 441448 626 441476 954
rect 442632 740 442684 746
rect 442632 682 442684 688
rect 441448 598 441568 626
rect 441540 480 441568 598
rect 442644 480 442672 682
rect 443748 610 443776 1294
rect 443840 746 443868 3060
rect 444944 1290 444972 3060
rect 445852 1352 445904 1358
rect 445852 1294 445904 1300
rect 444932 1284 444984 1290
rect 444932 1226 444984 1232
rect 445024 1216 445076 1222
rect 445024 1158 445076 1164
rect 443828 740 443880 746
rect 443828 682 443880 688
rect 443460 604 443512 610
rect 443460 546 443512 552
rect 443736 604 443788 610
rect 443736 546 443788 552
rect 437910 354 438022 480
rect 437584 326 438022 354
rect 437910 -960 438022 326
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443472 354 443500 546
rect 445036 480 445064 1158
rect 445760 1148 445812 1154
rect 445760 1090 445812 1096
rect 443798 354 443910 480
rect 443472 326 443910 354
rect 443798 -960 443910 326
rect 444994 -960 445106 480
rect 445772 270 445800 1090
rect 445864 354 445892 1294
rect 446048 1086 446076 3060
rect 446036 1080 446088 1086
rect 446036 1022 446088 1028
rect 447060 882 447088 3060
rect 447416 944 447468 950
rect 447416 886 447468 892
rect 447048 876 447100 882
rect 447048 818 447100 824
rect 447428 480 447456 886
rect 448256 678 448284 3060
rect 449360 1358 449388 3060
rect 449348 1352 449400 1358
rect 449348 1294 449400 1300
rect 450464 1222 450492 3060
rect 450452 1216 450504 1222
rect 450452 1158 450504 1164
rect 451568 1086 451596 3060
rect 451556 1080 451608 1086
rect 451556 1022 451608 1028
rect 448520 1012 448572 1018
rect 448704 1012 448756 1018
rect 448572 972 448704 1000
rect 448520 954 448572 960
rect 448704 954 448756 960
rect 451740 1012 451792 1018
rect 451740 954 451792 960
rect 450912 808 450964 814
rect 450912 750 450964 756
rect 448244 672 448296 678
rect 448244 614 448296 620
rect 449808 604 449860 610
rect 449808 546 449860 552
rect 449820 480 449848 546
rect 450924 480 450952 750
rect 446190 354 446302 480
rect 445864 326 446302 354
rect 445760 264 445812 270
rect 445760 206 445812 212
rect 446190 -960 446302 326
rect 447386 -960 447498 480
rect 448244 264 448296 270
rect 448582 218 448694 480
rect 448296 212 448694 218
rect 448244 206 448694 212
rect 448256 190 448694 206
rect 448582 -960 448694 190
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 451752 354 451780 954
rect 452078 354 452190 480
rect 451752 326 452190 354
rect 452078 -960 452190 326
rect 452580 202 452608 3060
rect 453212 1352 453264 1358
rect 453212 1294 453264 1300
rect 453224 1018 453252 1294
rect 453304 1148 453356 1154
rect 453304 1090 453356 1096
rect 453212 1012 453264 1018
rect 453212 954 453264 960
rect 453316 480 453344 1090
rect 452568 196 452620 202
rect 452568 138 452620 144
rect 453274 -960 453386 480
rect 453776 406 453804 3060
rect 454880 1290 454908 3060
rect 455696 1352 455748 1358
rect 455696 1294 455748 1300
rect 454868 1284 454920 1290
rect 454868 1226 454920 1232
rect 454132 740 454184 746
rect 454132 682 454184 688
rect 453764 400 453816 406
rect 453764 342 453816 348
rect 454144 354 454172 682
rect 455708 480 455736 1294
rect 455984 1154 456012 3060
rect 455972 1148 456024 1154
rect 455972 1090 456024 1096
rect 457088 1018 457116 3060
rect 457916 3046 458114 3074
rect 457076 1012 457128 1018
rect 457076 954 457128 960
rect 456892 944 456944 950
rect 456892 886 456944 892
rect 456904 480 456932 886
rect 454470 354 454582 480
rect 454144 326 454582 354
rect 454470 -960 454582 326
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 457916 338 457944 3046
rect 458088 876 458140 882
rect 458088 818 458140 824
rect 458100 480 458128 818
rect 459296 678 459324 3060
rect 460414 3046 460704 3074
rect 460020 944 460072 950
rect 460020 886 460072 892
rect 459192 672 459244 678
rect 459192 614 459244 620
rect 459284 672 459336 678
rect 459284 614 459336 620
rect 459204 480 459232 614
rect 457904 332 457956 338
rect 457904 274 457956 280
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460032 354 460060 886
rect 460358 354 460470 480
rect 460032 326 460470 354
rect 460358 -960 460470 326
rect 460676 134 460704 3046
rect 461504 610 461532 3060
rect 462608 1358 462636 3060
rect 462596 1352 462648 1358
rect 462596 1294 462648 1300
rect 461584 1216 461636 1222
rect 461584 1158 461636 1164
rect 461492 604 461544 610
rect 461492 546 461544 552
rect 461596 480 461624 1158
rect 462412 1080 462464 1086
rect 462412 1022 462464 1028
rect 460664 128 460716 134
rect 460664 70 460716 76
rect 461554 -960 461666 480
rect 462424 354 462452 1022
rect 462750 354 462862 480
rect 462424 326 462862 354
rect 462750 -960 462862 326
rect 463620 66 463648 3060
rect 463946 218 464058 480
rect 464816 474 464844 3060
rect 464804 468 464856 474
rect 464804 410 464856 416
rect 464988 400 465040 406
rect 465142 354 465254 480
rect 465040 348 465254 354
rect 464988 342 465254 348
rect 465000 326 465254 342
rect 463946 202 464200 218
rect 463946 196 464212 202
rect 463946 190 464160 196
rect 463608 60 463660 66
rect 463608 2 463660 8
rect 463946 -960 464058 190
rect 464160 138 464212 144
rect 465142 -960 465254 326
rect 465920 270 465948 3060
rect 466000 1284 466052 1290
rect 466000 1226 466052 1232
rect 466012 354 466040 1226
rect 466246 354 466358 480
rect 466012 326 466358 354
rect 465908 264 465960 270
rect 465908 206 465960 212
rect 466246 -960 466358 326
rect 467024 202 467052 3060
rect 467472 1148 467524 1154
rect 467472 1090 467524 1096
rect 467484 480 467512 1090
rect 468128 746 468156 3060
rect 469140 1290 469168 3060
rect 469128 1284 469180 1290
rect 469128 1226 469180 1232
rect 468300 1012 468352 1018
rect 468300 954 468352 960
rect 468116 740 468168 746
rect 468116 682 468168 688
rect 467012 196 467064 202
rect 467012 138 467064 144
rect 467442 -960 467554 480
rect 468312 354 468340 954
rect 470336 542 470364 3060
rect 471440 678 471468 3060
rect 471060 672 471112 678
rect 471060 614 471112 620
rect 471428 672 471480 678
rect 471428 614 471480 620
rect 470324 536 470376 542
rect 468638 354 468750 480
rect 468312 326 468750 354
rect 468638 -960 468750 326
rect 469834 354 469946 480
rect 470324 478 470376 484
rect 471072 480 471100 614
rect 469834 338 470088 354
rect 469834 332 470100 338
rect 469834 326 470048 332
rect 469834 -960 469946 326
rect 470048 274 470100 280
rect 471030 -960 471142 480
rect 472226 82 472338 480
rect 472544 406 472572 3060
rect 473452 604 473504 610
rect 473452 546 473504 552
rect 473464 480 473492 546
rect 472532 400 472584 406
rect 472532 342 472584 348
rect 472440 128 472492 134
rect 472226 76 472440 82
rect 472226 70 472492 76
rect 472226 54 472480 70
rect 472226 -960 472338 54
rect 473422 -960 473534 480
rect 473648 134 473676 3060
rect 474188 1352 474240 1358
rect 474188 1294 474240 1300
rect 474200 354 474228 1294
rect 474660 1154 474688 3060
rect 475856 1358 475884 3060
rect 476974 3046 477264 3074
rect 478078 3046 478368 3074
rect 475844 1352 475896 1358
rect 475844 1294 475896 1300
rect 474648 1148 474700 1154
rect 474648 1090 474700 1096
rect 474526 354 474638 480
rect 474200 326 474638 354
rect 473636 128 473688 134
rect 473636 70 473688 76
rect 474526 -960 474638 326
rect 475722 82 475834 480
rect 476580 468 476632 474
rect 476580 410 476632 416
rect 476592 354 476620 410
rect 476918 354 477030 480
rect 476592 326 477030 354
rect 475722 66 475976 82
rect 475722 60 475988 66
rect 475722 54 475936 60
rect 475722 -960 475834 54
rect 475936 2 475988 8
rect 476918 -960 477030 326
rect 477236 66 477264 3046
rect 478114 218 478226 480
rect 478340 474 478368 3046
rect 478328 468 478380 474
rect 478328 410 478380 416
rect 479168 338 479196 3060
rect 480180 678 480208 3060
rect 481390 3046 481588 3074
rect 481364 1284 481416 1290
rect 481364 1226 481416 1232
rect 480536 740 480588 746
rect 480536 682 480588 688
rect 479524 672 479576 678
rect 479524 614 479576 620
rect 480168 672 480220 678
rect 480168 614 480220 620
rect 479156 332 479208 338
rect 479156 274 479208 280
rect 478328 264 478380 270
rect 478114 212 478328 218
rect 479310 218 479422 480
rect 479536 406 479564 614
rect 480548 480 480576 682
rect 479524 400 479576 406
rect 479524 342 479576 348
rect 478114 206 478380 212
rect 478114 190 478368 206
rect 478984 202 479422 218
rect 478972 196 479422 202
rect 477224 60 477276 66
rect 477224 2 477276 8
rect 478114 -960 478226 190
rect 479024 190 479422 196
rect 478972 138 479024 144
rect 479310 -960 479422 190
rect 480506 -960 480618 480
rect 481376 354 481404 1226
rect 481560 950 481588 3046
rect 482480 1222 482508 3060
rect 482468 1216 482520 1222
rect 482468 1158 482520 1164
rect 481548 944 481600 950
rect 481548 886 481600 892
rect 483584 814 483612 3060
rect 483572 808 483624 814
rect 483572 750 483624 756
rect 482468 536 482520 542
rect 481702 354 481814 480
rect 482468 478 482520 484
rect 481376 326 481814 354
rect 482480 354 482508 478
rect 482806 354 482918 480
rect 482480 326 482918 354
rect 481702 -960 481814 326
rect 482806 -960 482918 326
rect 484002 354 484114 480
rect 484216 400 484268 406
rect 484002 348 484216 354
rect 484002 342 484268 348
rect 484002 326 484256 342
rect 484002 -960 484114 326
rect 484688 202 484716 3060
rect 485700 1086 485728 3060
rect 485688 1080 485740 1086
rect 485688 1022 485740 1028
rect 486896 1018 486924 3060
rect 488000 1154 488028 3060
rect 488816 1352 488868 1358
rect 488816 1294 488868 1300
rect 487252 1148 487304 1154
rect 487252 1090 487304 1096
rect 487988 1148 488040 1154
rect 487988 1090 488040 1096
rect 486884 1012 486936 1018
rect 486884 954 486936 960
rect 485198 354 485310 480
rect 484872 338 485310 354
rect 484860 332 485310 338
rect 484912 326 485310 332
rect 484860 274 484912 280
rect 484676 196 484728 202
rect 484676 138 484728 144
rect 485198 -960 485310 326
rect 486394 82 486506 480
rect 487264 354 487292 1090
rect 488828 480 488856 1294
rect 489104 746 489132 3060
rect 490208 1086 490236 3060
rect 490104 1080 490156 1086
rect 490104 1022 490156 1028
rect 490196 1080 490248 1086
rect 490196 1022 490248 1028
rect 489092 740 489144 746
rect 489092 682 489144 688
rect 490116 542 490144 1022
rect 491220 610 491248 3060
rect 492430 3046 492628 3074
rect 491208 604 491260 610
rect 491208 546 491260 552
rect 490104 536 490156 542
rect 487590 354 487702 480
rect 487264 326 487702 354
rect 486608 128 486660 134
rect 486394 76 486608 82
rect 486394 70 486660 76
rect 486394 54 486648 70
rect 486394 -960 486506 54
rect 487590 -960 487702 326
rect 488786 -960 488898 480
rect 489890 82 490002 480
rect 490104 478 490156 484
rect 490748 468 490800 474
rect 490748 410 490800 416
rect 490760 354 490788 410
rect 491086 354 491198 480
rect 490760 326 491198 354
rect 489890 66 490144 82
rect 489890 60 490156 66
rect 489890 54 490104 60
rect 489890 -960 490002 54
rect 490104 2 490156 8
rect 491086 -960 491198 326
rect 492282 218 492394 480
rect 492600 270 492628 3046
rect 493520 1358 493548 3060
rect 493508 1352 493560 1358
rect 493508 1294 493560 1300
rect 494624 950 494652 3060
rect 495728 1290 495756 3060
rect 495716 1284 495768 1290
rect 495716 1226 495768 1232
rect 495532 1216 495584 1222
rect 495532 1158 495584 1164
rect 494796 1080 494848 1086
rect 494796 1022 494848 1028
rect 494612 944 494664 950
rect 494612 886 494664 892
rect 494808 882 494836 1022
rect 494704 876 494756 882
rect 494704 818 494756 824
rect 494796 876 494848 882
rect 494796 818 494848 824
rect 493140 672 493192 678
rect 493140 614 493192 620
rect 493152 354 493180 614
rect 494716 480 494744 818
rect 493478 354 493590 480
rect 493152 326 493590 354
rect 492496 264 492548 270
rect 492282 212 492496 218
rect 492282 206 492548 212
rect 492588 264 492640 270
rect 492588 206 492640 212
rect 492282 190 492536 206
rect 492282 -960 492394 190
rect 493478 -960 493590 326
rect 494674 -960 494786 480
rect 495544 354 495572 1158
rect 495870 354 495982 480
rect 495544 326 495982 354
rect 495870 -960 495982 326
rect 496740 66 496768 3060
rect 497096 808 497148 814
rect 497096 750 497148 756
rect 497108 480 497136 750
rect 496728 60 496780 66
rect 496728 2 496780 8
rect 497066 -960 497178 480
rect 497936 474 497964 3060
rect 497924 468 497976 474
rect 497924 410 497976 416
rect 498170 218 498282 480
rect 499040 406 499068 3060
rect 499120 536 499172 542
rect 499120 478 499172 484
rect 499028 400 499080 406
rect 499028 342 499080 348
rect 499132 354 499160 478
rect 499366 354 499478 480
rect 499132 326 499478 354
rect 498170 202 498424 218
rect 498170 196 498436 202
rect 498170 190 498384 196
rect 498170 -960 498282 190
rect 498384 138 498436 144
rect 499366 -960 499478 326
rect 500144 134 500172 3060
rect 501248 1018 501276 3060
rect 501420 1148 501472 1154
rect 501420 1090 501472 1096
rect 500592 1012 500644 1018
rect 500592 954 500644 960
rect 501236 1012 501288 1018
rect 501236 954 501288 960
rect 500604 480 500632 954
rect 500132 128 500184 134
rect 500132 70 500184 76
rect 500562 -960 500674 480
rect 501432 354 501460 1090
rect 502260 678 502288 3060
rect 502984 740 503036 746
rect 502984 682 503036 688
rect 502248 672 502300 678
rect 502248 614 502300 620
rect 502996 480 503024 682
rect 503456 542 503484 3060
rect 503812 876 503864 882
rect 503812 818 503864 824
rect 503444 536 503496 542
rect 501758 354 501870 480
rect 501432 326 501870 354
rect 501758 -960 501870 326
rect 502954 -960 503066 480
rect 503444 478 503496 484
rect 503824 354 503852 818
rect 504150 354 504262 480
rect 503824 326 504262 354
rect 504560 338 504588 3060
rect 505376 604 505428 610
rect 505376 546 505428 552
rect 505388 480 505416 546
rect 504150 -960 504262 326
rect 504548 332 504600 338
rect 504548 274 504600 280
rect 505346 -960 505458 480
rect 505664 202 505692 3060
rect 506768 1222 506796 3060
rect 507308 1352 507360 1358
rect 507308 1294 507360 1300
rect 506756 1216 506808 1222
rect 506756 1158 506808 1164
rect 506450 218 506562 480
rect 507320 354 507348 1294
rect 507780 1154 507808 3060
rect 507768 1148 507820 1154
rect 507768 1090 507820 1096
rect 508872 944 508924 950
rect 508872 886 508924 892
rect 508884 480 508912 886
rect 508976 610 509004 3060
rect 510080 1290 510108 3060
rect 511198 3046 511488 3074
rect 512302 3046 512684 3074
rect 513406 3058 513512 3074
rect 532608 3062 532660 3068
rect 540796 3120 540848 3126
rect 540796 3062 540848 3068
rect 513406 3052 513524 3058
rect 513406 3046 513472 3052
rect 509700 1284 509752 1290
rect 509700 1226 509752 1232
rect 510068 1284 510120 1290
rect 510068 1226 510120 1232
rect 508964 604 509016 610
rect 508964 546 509016 552
rect 507646 354 507758 480
rect 507320 326 507758 354
rect 506664 264 506716 270
rect 506450 212 506664 218
rect 506450 206 506716 212
rect 505652 196 505704 202
rect 505652 138 505704 144
rect 506450 190 506704 206
rect 506450 -960 506562 190
rect 507646 -960 507758 326
rect 508842 -960 508954 480
rect 509712 354 509740 1226
rect 510038 354 510150 480
rect 509712 326 510150 354
rect 510038 -960 510150 326
rect 511234 82 511346 480
rect 511460 270 511488 3046
rect 512092 468 512144 474
rect 512092 410 512144 416
rect 512104 354 512132 410
rect 512430 354 512542 480
rect 512104 326 512542 354
rect 511448 264 511500 270
rect 511448 206 511500 212
rect 511234 66 511488 82
rect 511234 60 511500 66
rect 511234 54 511448 60
rect 511234 -960 511346 54
rect 511448 2 511500 8
rect 512430 -960 512542 326
rect 512656 66 512684 3046
rect 513472 2994 513524 3000
rect 514496 814 514524 3060
rect 514852 2984 514904 2990
rect 514852 2926 514904 2932
rect 514760 2916 514812 2922
rect 514760 2858 514812 2864
rect 514772 1154 514800 2858
rect 514864 1222 514892 2926
rect 514852 1216 514904 1222
rect 514852 1158 514904 1164
rect 514760 1148 514812 1154
rect 514760 1090 514812 1096
rect 515600 1018 515628 3060
rect 515496 1012 515548 1018
rect 515496 954 515548 960
rect 515588 1012 515640 1018
rect 515588 954 515640 960
rect 514484 808 514536 814
rect 514484 750 514536 756
rect 513380 400 513432 406
rect 513534 354 513646 480
rect 513432 348 513646 354
rect 513380 342 513646 348
rect 513392 326 513646 342
rect 512644 60 512696 66
rect 512644 2 512696 8
rect 513534 -960 513646 326
rect 514730 82 514842 480
rect 515508 354 515536 954
rect 515926 354 516038 480
rect 516704 474 516732 3060
rect 517152 672 517204 678
rect 517152 614 517204 620
rect 517164 480 517192 614
rect 516692 468 516744 474
rect 516692 410 516744 416
rect 515508 326 516038 354
rect 514944 128 514996 134
rect 514730 76 514944 82
rect 514730 70 514996 76
rect 514730 54 514984 70
rect 514730 -960 514842 54
rect 515926 -960 516038 326
rect 517122 -960 517234 480
rect 517808 406 517836 3060
rect 517980 536 518032 542
rect 517980 478 518032 484
rect 517796 400 517848 406
rect 517796 342 517848 348
rect 517992 354 518020 478
rect 518318 354 518430 480
rect 517992 326 518430 354
rect 518318 -960 518430 326
rect 518820 134 518848 3060
rect 520016 950 520044 3060
rect 520188 2848 520240 2854
rect 520188 2790 520240 2796
rect 520200 1290 520228 2790
rect 520188 1284 520240 1290
rect 520188 1226 520240 1232
rect 520004 944 520056 950
rect 520004 886 520056 892
rect 519514 354 519626 480
rect 519514 338 519768 354
rect 519514 332 519780 338
rect 519514 326 519728 332
rect 518808 128 518860 134
rect 518808 70 518860 76
rect 519514 -960 519626 326
rect 519728 274 519780 280
rect 520710 218 520822 480
rect 521120 338 521148 3060
rect 521844 2984 521896 2990
rect 521844 2926 521896 2932
rect 521856 480 521884 2926
rect 522224 746 522252 3060
rect 523040 2916 523092 2922
rect 523040 2858 523092 2864
rect 522212 740 522264 746
rect 522212 682 522264 688
rect 523052 480 523080 2858
rect 523328 882 523356 3060
rect 524340 1290 524368 3060
rect 525432 2780 525484 2786
rect 525432 2722 525484 2728
rect 524328 1284 524380 1290
rect 524328 1226 524380 1232
rect 523316 876 523368 882
rect 523316 818 523368 824
rect 524236 604 524288 610
rect 524236 546 524288 552
rect 524248 480 524276 546
rect 525444 480 525472 2722
rect 525536 1086 525564 3060
rect 525800 2916 525852 2922
rect 525800 2858 525852 2864
rect 525524 1080 525576 1086
rect 525524 1022 525576 1028
rect 525812 1018 525840 2858
rect 526640 1358 526668 3060
rect 526628 1352 526680 1358
rect 526628 1294 526680 1300
rect 527744 1018 527772 3060
rect 528848 1222 528876 3060
rect 529020 3052 529072 3058
rect 529020 2994 529072 3000
rect 528836 1216 528888 1222
rect 528836 1158 528888 1164
rect 525800 1012 525852 1018
rect 525800 954 525852 960
rect 527732 1012 527784 1018
rect 527732 954 527784 960
rect 529032 480 529060 2994
rect 529756 808 529808 814
rect 529756 750 529808 756
rect 521108 332 521160 338
rect 521108 274 521160 280
rect 520384 202 520822 218
rect 520372 196 520822 202
rect 520424 190 520822 196
rect 520372 138 520424 144
rect 520710 -960 520822 190
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526260 264 526312 270
rect 526598 218 526710 480
rect 526312 212 526710 218
rect 526260 206 526710 212
rect 526272 190 526710 206
rect 526598 -960 526710 190
rect 527794 82 527906 480
rect 527794 66 528048 82
rect 527794 60 528060 66
rect 527794 54 528008 60
rect 527794 -960 527906 54
rect 528008 2 528060 8
rect 528990 -960 529102 480
rect 529768 354 529796 750
rect 530094 354 530206 480
rect 529768 326 530206 354
rect 530094 -960 530206 326
rect 531056 66 531084 3060
rect 531320 2916 531372 2922
rect 531320 2858 531372 2864
rect 531332 480 531360 2858
rect 532160 814 532188 3060
rect 532240 2916 532292 2922
rect 532240 2858 532292 2864
rect 532252 882 532280 2858
rect 532620 1290 532648 3062
rect 532608 1284 532660 1290
rect 532608 1226 532660 1232
rect 533264 1154 533292 3060
rect 533252 1148 533304 1154
rect 533252 1090 533304 1096
rect 532240 876 532292 882
rect 532240 818 532292 824
rect 532148 808 532200 814
rect 532148 750 532200 756
rect 531044 60 531096 66
rect 531044 2 531096 8
rect 531290 -960 531402 480
rect 532148 468 532200 474
rect 532148 410 532200 416
rect 532160 354 532188 410
rect 532486 354 532598 480
rect 532160 326 532598 354
rect 532486 -960 532598 326
rect 533682 354 533794 480
rect 534368 406 534396 3060
rect 533896 400 533948 406
rect 533682 348 533896 354
rect 533682 342 533948 348
rect 534356 400 534408 406
rect 534356 342 534408 348
rect 533682 326 533936 342
rect 533682 -960 533794 326
rect 534540 128 534592 134
rect 534878 82 534990 480
rect 535380 270 535408 3060
rect 535552 3052 535604 3058
rect 535552 2994 535604 3000
rect 535564 1358 535592 2994
rect 536576 2990 536604 3060
rect 536564 2984 536616 2990
rect 536564 2926 536616 2932
rect 536840 2848 536892 2854
rect 536840 2790 536892 2796
rect 535552 1352 535604 1358
rect 535552 1294 535604 1300
rect 536852 1086 536880 2790
rect 536840 1080 536892 1086
rect 536840 1022 536892 1028
rect 536104 944 536156 950
rect 536104 886 536156 892
rect 536116 480 536144 886
rect 535368 264 535420 270
rect 535368 206 535420 212
rect 534592 76 534990 82
rect 534540 70 534990 76
rect 534552 54 534990 70
rect 534878 -960 534990 54
rect 536074 -960 536186 480
rect 537178 354 537290 480
rect 537178 338 537432 354
rect 537178 332 537444 338
rect 537178 326 537392 332
rect 537178 -960 537290 326
rect 537392 274 537444 280
rect 537680 202 537708 3060
rect 538220 740 538272 746
rect 538220 682 538272 688
rect 538232 354 538260 682
rect 538374 354 538486 480
rect 538232 326 538486 354
rect 538784 338 538812 3060
rect 539600 2916 539652 2922
rect 539600 2858 539652 2864
rect 539612 480 539640 2858
rect 539888 1358 539916 3060
rect 539876 1352 539928 1358
rect 539876 1294 539928 1300
rect 540808 480 540836 3062
rect 540900 746 540928 3060
rect 541992 2916 542044 2922
rect 541992 2858 542044 2864
rect 541532 2848 541584 2854
rect 541532 2790 541584 2796
rect 541544 1154 541572 2790
rect 541532 1148 541584 1154
rect 541532 1090 541584 1096
rect 540888 740 540940 746
rect 540888 682 540940 688
rect 542004 480 542032 2858
rect 542096 678 542124 3060
rect 543214 3058 543504 3074
rect 542820 3052 542872 3058
rect 543214 3052 543516 3058
rect 543214 3046 543464 3052
rect 542820 2994 542872 3000
rect 544318 3046 544608 3074
rect 543464 2994 543516 3000
rect 542084 672 542136 678
rect 542084 614 542136 620
rect 537668 196 537720 202
rect 537668 138 537720 144
rect 538374 -960 538486 326
rect 538772 332 538824 338
rect 538772 274 538824 280
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 542832 354 542860 2994
rect 544384 1012 544436 1018
rect 544384 954 544436 960
rect 544396 480 544424 954
rect 544580 542 544608 3046
rect 545408 610 545436 3060
rect 545488 1216 545540 1222
rect 545488 1158 545540 1164
rect 545396 604 545448 610
rect 545396 546 545448 552
rect 544568 536 544620 542
rect 543158 354 543270 480
rect 542832 326 543270 354
rect 543158 -960 543270 326
rect 544354 -960 544466 480
rect 544568 478 544620 484
rect 545500 480 545528 1158
rect 545458 -960 545570 480
rect 546420 134 546448 3060
rect 546696 480 546724 3198
rect 556462 3182 556752 3198
rect 560878 3194 561168 3210
rect 560878 3188 561180 3194
rect 560878 3182 561128 3188
rect 561128 3130 561180 3136
rect 563152 3120 563204 3126
rect 547616 882 547644 3060
rect 548734 3046 548932 3074
rect 547604 876 547656 882
rect 547604 818 547656 824
rect 548708 808 548760 814
rect 548708 750 548760 756
rect 546408 128 546460 134
rect 546408 70 546460 76
rect 546654 -960 546766 480
rect 547850 82 547962 480
rect 548720 354 548748 750
rect 548904 474 548932 3046
rect 550272 2848 550324 2854
rect 550272 2790 550324 2796
rect 550284 480 550312 2790
rect 550928 814 550956 3060
rect 550916 808 550968 814
rect 550916 750 550968 756
rect 548892 468 548944 474
rect 548892 410 548944 416
rect 549046 354 549158 480
rect 548720 326 549158 354
rect 547850 66 548104 82
rect 547850 60 548116 66
rect 547850 54 548064 60
rect 547850 -960 547962 54
rect 548064 2 548116 8
rect 549046 -960 549158 326
rect 550242 -960 550354 480
rect 551100 400 551152 406
rect 551438 354 551550 480
rect 551152 348 551550 354
rect 551100 342 551550 348
rect 551112 326 551550 342
rect 551438 -960 551550 326
rect 551940 66 551968 3060
rect 553768 2984 553820 2990
rect 553768 2926 553820 2932
rect 553780 480 553808 2926
rect 552634 218 552746 480
rect 552848 264 552900 270
rect 552634 212 552848 218
rect 552634 206 552900 212
rect 552634 190 552888 206
rect 551928 60 551980 66
rect 551928 2 551980 8
rect 552634 -960 552746 190
rect 553738 -960 553850 480
rect 554240 270 554268 3060
rect 554228 264 554280 270
rect 554934 218 555046 480
rect 555344 406 555372 3060
rect 557184 3046 557474 3074
rect 558670 3046 558868 3074
rect 563086 3068 563152 3074
rect 563086 3062 563204 3068
rect 556988 1352 557040 1358
rect 556988 1294 557040 1300
rect 555332 400 555384 406
rect 555332 342 555384 348
rect 556130 354 556242 480
rect 554228 206 554280 212
rect 554792 202 555046 218
rect 554780 196 555046 202
rect 554832 190 555046 196
rect 554780 138 554832 144
rect 554934 -960 555046 190
rect 556130 338 556384 354
rect 556130 332 556396 338
rect 556130 326 556344 332
rect 556130 -960 556242 326
rect 556344 274 556396 280
rect 557000 218 557028 1294
rect 557184 338 557212 3046
rect 558552 740 558604 746
rect 558552 682 558604 688
rect 558564 480 558592 682
rect 557172 332 557224 338
rect 557172 274 557224 280
rect 557326 218 557438 480
rect 557000 190 557438 218
rect 557326 -960 557438 190
rect 558522 -960 558634 480
rect 558840 202 558868 3046
rect 559760 2854 559788 3060
rect 560484 3052 560536 3058
rect 560484 2994 560536 3000
rect 559748 2848 559800 2854
rect 559748 2790 559800 2796
rect 559748 672 559800 678
rect 559748 614 559800 620
rect 559760 480 559788 614
rect 558828 196 558880 202
rect 558828 138 558880 144
rect 559718 -960 559830 480
rect 560496 354 560524 2994
rect 561968 2922 561996 3060
rect 563086 3046 563192 3062
rect 564190 3058 564388 3074
rect 564190 3052 564400 3058
rect 564190 3046 564348 3052
rect 564348 2994 564400 3000
rect 561956 2916 562008 2922
rect 561956 2858 562008 2864
rect 565636 876 565688 882
rect 565636 818 565688 824
rect 563244 672 563296 678
rect 563244 614 563296 620
rect 562048 604 562100 610
rect 562048 546 562100 552
rect 562060 480 562088 546
rect 563256 480 563284 614
rect 565648 480 565676 818
rect 568040 480 568068 3266
rect 569132 808 569184 814
rect 569132 750 569184 756
rect 569144 480 569172 750
rect 571536 480 571564 3334
rect 575112 3256 575164 3262
rect 575112 3198 575164 3204
rect 575124 480 575152 3198
rect 579804 3188 579856 3194
rect 579804 3130 579856 3136
rect 578608 2848 578660 2854
rect 578608 2790 578660 2796
rect 578620 480 578648 2790
rect 579816 480 579844 3130
rect 582196 3120 582248 3126
rect 582196 3062 582248 3068
rect 581000 2916 581052 2922
rect 581000 2858 581052 2864
rect 581012 480 581040 2858
rect 582208 480 582236 3062
rect 583392 3052 583444 3058
rect 583392 2994 583444 3000
rect 583404 480 583432 2994
rect 560822 354 560934 480
rect 560496 326 560934 354
rect 560822 -960 560934 326
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 82 564522 480
rect 564624 128 564676 134
rect 564410 76 564624 82
rect 564410 70 564676 76
rect 564410 54 564664 70
rect 564410 -960 564522 54
rect 565606 -960 565718 480
rect 566802 354 566914 480
rect 567016 468 567068 474
rect 567016 410 567068 416
rect 567028 354 567056 410
rect 566802 326 567056 354
rect 566802 -960 566914 326
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 82 570410 480
rect 570298 66 570552 82
rect 570298 60 570564 66
rect 570298 54 570512 60
rect 570298 -960 570410 54
rect 570512 2 570564 8
rect 571494 -960 571606 480
rect 572690 218 572802 480
rect 573548 400 573600 406
rect 573886 354 573998 480
rect 573600 348 573998 354
rect 573548 342 573998 348
rect 573560 326 573998 342
rect 572904 264 572956 270
rect 572690 212 572904 218
rect 572690 206 572956 212
rect 572690 190 572944 206
rect 572690 -960 572802 190
rect 573886 -960 573998 326
rect 575082 -960 575194 480
rect 576278 354 576390 480
rect 575952 338 576390 354
rect 575940 332 576390 338
rect 575992 326 576390 332
rect 575940 274 575992 280
rect 576278 -960 576390 326
rect 577382 218 577494 480
rect 577148 202 577494 218
rect 577136 196 577494 202
rect 577188 190 577494 196
rect 577136 138 577188 144
rect 577382 -960 577494 190
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 2778 697312 2834 697368
rect 581642 697176 581698 697232
rect 581642 691464 581698 691520
rect 2778 690784 2834 690840
rect 2778 684256 2834 684312
rect 582378 683848 582434 683904
rect 582378 678408 582434 678464
rect 2778 678000 2834 678056
rect 2778 671200 2834 671256
rect 582378 670656 582434 670712
rect 582378 665352 582434 665408
rect 2778 665216 2834 665272
rect 2778 658144 2834 658200
rect 582378 657328 582434 657384
rect 2778 652432 2834 652488
rect 582378 652296 582434 652352
rect 2778 645088 2834 645144
rect 581642 644000 581698 644056
rect 2778 639648 2834 639704
rect 581642 639240 581698 639296
rect 2778 632032 2834 632088
rect 582378 630808 582434 630864
rect 2778 626864 2834 626920
rect 582378 626184 582434 626240
rect 2778 619112 2834 619168
rect 581642 617480 581698 617536
rect 2778 613944 2834 614000
rect 581642 613128 581698 613184
rect 2778 606056 2834 606112
rect 581642 604152 581698 604208
rect 2778 601296 2834 601352
rect 581642 600072 581698 600128
rect 1582 593000 1638 593056
rect 581642 590960 581698 591016
rect 1582 588512 1638 588568
rect 581642 587016 581698 587072
rect 2042 579944 2098 580000
rect 581642 577632 581698 577688
rect 2042 575728 2098 575784
rect 581642 573960 581698 574016
rect 1490 566888 1546 566944
rect 582378 564304 582434 564360
rect 1490 562944 1546 563000
rect 582378 560904 582434 560960
rect 1490 553832 1546 553888
rect 581642 551112 581698 551168
rect 1490 550160 1546 550216
rect 581642 547712 581698 547768
rect 1398 540776 1454 540832
rect 582378 537784 582434 537840
rect 1398 537376 1454 537432
rect 582378 534792 582434 534848
rect 1490 527856 1546 527912
rect 1490 524592 1546 524648
rect 582378 524456 582434 524512
rect 582378 521736 582434 521792
rect 1582 514800 1638 514856
rect 1582 511808 1638 511864
rect 582378 511264 582434 511320
rect 582378 508680 582434 508736
rect 1582 501744 1638 501800
rect 1582 499024 1638 499080
rect 581642 497936 581698 497992
rect 581642 495624 581698 495680
rect 1582 488688 1638 488744
rect 1582 486240 1638 486296
rect 582378 484608 582434 484664
rect 582378 482568 582434 482624
rect 2778 475632 2834 475688
rect 2778 473456 2834 473512
rect 581642 471416 581698 471472
rect 581642 469512 581698 469568
rect 1582 462576 1638 462632
rect 1582 460672 1638 460728
rect 581642 458088 581698 458144
rect 581642 456456 581698 456512
rect 2778 449520 2834 449576
rect 2778 447888 2834 447944
rect 2778 436600 2834 436656
rect 2778 435104 2834 435160
rect 2778 423544 2834 423600
rect 2778 422320 2834 422376
rect 1306 294344 1362 294400
rect 1306 293120 1362 293176
rect 2778 281560 2834 281616
rect 2778 280064 2834 280120
rect 1306 268776 1362 268832
rect 1306 267144 1362 267200
rect 582378 260480 582434 260536
rect 582378 258848 582434 258904
rect 1306 255992 1362 256048
rect 1306 254088 1362 254144
rect 580906 247016 580962 247072
rect 580906 245520 580962 245576
rect 2778 243208 2834 243264
rect 2778 241032 2834 241088
rect 582378 234368 582434 234424
rect 582378 232328 582434 232384
rect 2778 230560 2834 230616
rect 2778 227976 2834 228032
rect 580906 220904 580962 220960
rect 580906 219000 580962 219056
rect 2778 217640 2834 217696
rect 2778 214920 2834 214976
rect 582378 208256 582434 208312
rect 582378 205672 582434 205728
rect 2778 204856 2834 204912
rect 2778 201864 2834 201920
rect 580906 194656 580962 194712
rect 580906 192480 580962 192536
rect 1306 192072 1362 192128
rect 1306 188808 1362 188864
rect 580906 182416 580962 182472
rect 2778 179288 2834 179344
rect 580906 179152 580962 179208
rect 2778 175888 2834 175944
rect 580906 168544 580962 168600
rect 2778 166504 2834 166560
rect 580906 165824 580962 165880
rect 2778 162832 2834 162888
rect 580906 156304 580962 156360
rect 1306 153720 1362 153776
rect 580906 152632 580962 152688
rect 1306 149776 1362 149832
rect 580906 142568 580962 142624
rect 570 140936 626 140992
rect 580906 139304 580962 139360
rect 570 136720 626 136776
rect 580906 130192 580962 130248
rect 754 128152 810 128208
rect 580906 125976 580962 126032
rect 754 123664 810 123720
rect 579894 116320 579950 116376
rect 1306 115368 1362 115424
rect 579894 112784 579950 112840
rect 1306 110608 1362 110664
rect 580906 103536 580962 103592
rect 1582 102584 1638 102640
rect 580906 99456 580962 99512
rect 1582 97552 1638 97608
rect 580906 90208 580962 90264
rect 1582 89800 1638 89856
rect 580906 86128 580962 86184
rect 1582 84632 1638 84688
rect 579894 77288 579950 77344
rect 1582 77016 1638 77072
rect 579894 72936 579950 72992
rect 1582 71576 1638 71632
rect 1490 64232 1546 64288
rect 580906 64096 580962 64152
rect 580906 59608 580962 59664
rect 1490 58520 1546 58576
rect 2042 51448 2098 51504
rect 580906 51040 580962 51096
rect 580906 46280 580962 46336
rect 2042 45464 2098 45520
rect 2042 38664 2098 38720
rect 580906 37984 580962 38040
rect 580906 33088 580962 33144
rect 2042 32408 2098 32464
rect 1490 25880 1546 25936
rect 580906 24928 580962 24984
rect 580906 19760 580962 19816
rect 1490 19352 1546 19408
rect 2042 13096 2098 13152
rect 582378 12416 582434 12472
rect 582378 6568 582434 6624
rect 2042 6432 2098 6488
rect 6274 176 6330 232
rect 5446 40 5502 96
rect 12162 448 12218 504
rect 13726 312 13782 368
rect 23938 40 23994 96
rect 25042 176 25098 232
rect 25686 176 25742 232
rect 28906 584 28962 640
rect 30838 448 30894 504
rect 31942 312 31998 368
rect 37002 40 37058 96
rect 42706 176 42762 232
rect 46294 584 46350 640
rect 46846 176 46902 232
rect 54022 40 54078 96
rect 62854 176 62910 232
<< metal3 >>
rect -960 697370 480 697460
rect 2773 697370 2839 697373
rect -960 697368 2839 697370
rect -960 697312 2778 697368
rect 2834 697312 2839 697368
rect -960 697310 2839 697312
rect -960 697220 480 697310
rect 2773 697307 2839 697310
rect 581637 697234 581703 697237
rect 583520 697234 584960 697324
rect 581637 697232 584960 697234
rect 581637 697176 581642 697232
rect 581698 697176 584960 697232
rect 581637 697174 584960 697176
rect 581637 697171 581703 697174
rect 583520 697084 584960 697174
rect 581637 691522 581703 691525
rect 580796 691520 581703 691522
rect 580796 691464 581642 691520
rect 581698 691464 581703 691520
rect 580796 691462 581703 691464
rect 581637 691459 581703 691462
rect 2773 690842 2839 690845
rect 2773 690840 3220 690842
rect 2773 690784 2778 690840
rect 2834 690784 3220 690840
rect 2773 690782 3220 690784
rect 2773 690779 2839 690782
rect -960 684314 480 684404
rect 2773 684314 2839 684317
rect -960 684312 2839 684314
rect -960 684256 2778 684312
rect 2834 684256 2839 684312
rect -960 684254 2839 684256
rect -960 684164 480 684254
rect 2773 684251 2839 684254
rect 582373 683906 582439 683909
rect 583520 683906 584960 683996
rect 582373 683904 584960 683906
rect 582373 683848 582378 683904
rect 582434 683848 584960 683904
rect 582373 683846 584960 683848
rect 582373 683843 582439 683846
rect 583520 683756 584960 683846
rect 582373 678466 582439 678469
rect 580796 678464 582439 678466
rect 580796 678408 582378 678464
rect 582434 678408 582439 678464
rect 580796 678406 582439 678408
rect 582373 678403 582439 678406
rect 2773 678058 2839 678061
rect 2773 678056 3220 678058
rect 2773 678000 2778 678056
rect 2834 678000 3220 678056
rect 2773 677998 3220 678000
rect 2773 677995 2839 677998
rect -960 671258 480 671348
rect 2773 671258 2839 671261
rect -960 671256 2839 671258
rect -960 671200 2778 671256
rect 2834 671200 2839 671256
rect -960 671198 2839 671200
rect -960 671108 480 671198
rect 2773 671195 2839 671198
rect 582373 670714 582439 670717
rect 583520 670714 584960 670804
rect 582373 670712 584960 670714
rect 582373 670656 582378 670712
rect 582434 670656 584960 670712
rect 582373 670654 584960 670656
rect 582373 670651 582439 670654
rect 583520 670564 584960 670654
rect 582373 665410 582439 665413
rect 580796 665408 582439 665410
rect 580796 665352 582378 665408
rect 582434 665352 582439 665408
rect 580796 665350 582439 665352
rect 582373 665347 582439 665350
rect 2773 665274 2839 665277
rect 2773 665272 3220 665274
rect 2773 665216 2778 665272
rect 2834 665216 3220 665272
rect 2773 665214 3220 665216
rect 2773 665211 2839 665214
rect -960 658202 480 658292
rect 2773 658202 2839 658205
rect -960 658200 2839 658202
rect -960 658144 2778 658200
rect 2834 658144 2839 658200
rect -960 658142 2839 658144
rect -960 658052 480 658142
rect 2773 658139 2839 658142
rect 582373 657386 582439 657389
rect 583520 657386 584960 657476
rect 582373 657384 584960 657386
rect 582373 657328 582378 657384
rect 582434 657328 584960 657384
rect 582373 657326 584960 657328
rect 582373 657323 582439 657326
rect 583520 657236 584960 657326
rect 2773 652490 2839 652493
rect 2773 652488 3220 652490
rect 2773 652432 2778 652488
rect 2834 652432 3220 652488
rect 2773 652430 3220 652432
rect 2773 652427 2839 652430
rect 582373 652354 582439 652357
rect 580796 652352 582439 652354
rect 580796 652296 582378 652352
rect 582434 652296 582439 652352
rect 580796 652294 582439 652296
rect 582373 652291 582439 652294
rect -960 645146 480 645236
rect 2773 645146 2839 645149
rect -960 645144 2839 645146
rect -960 645088 2778 645144
rect 2834 645088 2839 645144
rect -960 645086 2839 645088
rect -960 644996 480 645086
rect 2773 645083 2839 645086
rect 581637 644058 581703 644061
rect 583520 644058 584960 644148
rect 581637 644056 584960 644058
rect 581637 644000 581642 644056
rect 581698 644000 584960 644056
rect 581637 643998 584960 644000
rect 581637 643995 581703 643998
rect 583520 643908 584960 643998
rect 2773 639706 2839 639709
rect 2773 639704 3220 639706
rect 2773 639648 2778 639704
rect 2834 639648 3220 639704
rect 2773 639646 3220 639648
rect 2773 639643 2839 639646
rect 581637 639298 581703 639301
rect 580796 639296 581703 639298
rect 580796 639240 581642 639296
rect 581698 639240 581703 639296
rect 580796 639238 581703 639240
rect 581637 639235 581703 639238
rect -960 632090 480 632180
rect 2773 632090 2839 632093
rect -960 632088 2839 632090
rect -960 632032 2778 632088
rect 2834 632032 2839 632088
rect -960 632030 2839 632032
rect -960 631940 480 632030
rect 2773 632027 2839 632030
rect 582373 630866 582439 630869
rect 583520 630866 584960 630956
rect 582373 630864 584960 630866
rect 582373 630808 582378 630864
rect 582434 630808 584960 630864
rect 582373 630806 584960 630808
rect 582373 630803 582439 630806
rect 583520 630716 584960 630806
rect 2773 626922 2839 626925
rect 2773 626920 3220 626922
rect 2773 626864 2778 626920
rect 2834 626864 3220 626920
rect 2773 626862 3220 626864
rect 2773 626859 2839 626862
rect 582373 626242 582439 626245
rect 580796 626240 582439 626242
rect 580796 626184 582378 626240
rect 582434 626184 582439 626240
rect 580796 626182 582439 626184
rect 582373 626179 582439 626182
rect -960 619170 480 619260
rect 2773 619170 2839 619173
rect -960 619168 2839 619170
rect -960 619112 2778 619168
rect 2834 619112 2839 619168
rect -960 619110 2839 619112
rect -960 619020 480 619110
rect 2773 619107 2839 619110
rect 581637 617538 581703 617541
rect 583520 617538 584960 617628
rect 581637 617536 584960 617538
rect 581637 617480 581642 617536
rect 581698 617480 584960 617536
rect 581637 617478 584960 617480
rect 581637 617475 581703 617478
rect 583520 617388 584960 617478
rect 2773 614002 2839 614005
rect 2773 614000 3220 614002
rect 2773 613944 2778 614000
rect 2834 613944 3220 614000
rect 2773 613942 3220 613944
rect 2773 613939 2839 613942
rect 581637 613186 581703 613189
rect 580796 613184 581703 613186
rect 580796 613128 581642 613184
rect 581698 613128 581703 613184
rect 580796 613126 581703 613128
rect 581637 613123 581703 613126
rect -960 606114 480 606204
rect 2773 606114 2839 606117
rect -960 606112 2839 606114
rect -960 606056 2778 606112
rect 2834 606056 2839 606112
rect -960 606054 2839 606056
rect -960 605964 480 606054
rect 2773 606051 2839 606054
rect 581637 604210 581703 604213
rect 583520 604210 584960 604300
rect 581637 604208 584960 604210
rect 581637 604152 581642 604208
rect 581698 604152 584960 604208
rect 581637 604150 584960 604152
rect 581637 604147 581703 604150
rect 583520 604060 584960 604150
rect 2773 601354 2839 601357
rect 2773 601352 3220 601354
rect 2773 601296 2778 601352
rect 2834 601296 3220 601352
rect 2773 601294 3220 601296
rect 2773 601291 2839 601294
rect 581637 600130 581703 600133
rect 580796 600128 581703 600130
rect 580796 600072 581642 600128
rect 581698 600072 581703 600128
rect 580796 600070 581703 600072
rect 581637 600067 581703 600070
rect -960 593058 480 593148
rect 1577 593058 1643 593061
rect -960 593056 1643 593058
rect -960 593000 1582 593056
rect 1638 593000 1643 593056
rect -960 592998 1643 593000
rect -960 592908 480 592998
rect 1577 592995 1643 592998
rect 581637 591018 581703 591021
rect 583520 591018 584960 591108
rect 581637 591016 584960 591018
rect 581637 590960 581642 591016
rect 581698 590960 584960 591016
rect 581637 590958 584960 590960
rect 581637 590955 581703 590958
rect 583520 590868 584960 590958
rect 1577 588570 1643 588573
rect 1577 588568 3220 588570
rect 1577 588512 1582 588568
rect 1638 588512 3220 588568
rect 1577 588510 3220 588512
rect 1577 588507 1643 588510
rect 581637 587074 581703 587077
rect 580796 587072 581703 587074
rect 580796 587016 581642 587072
rect 581698 587016 581703 587072
rect 580796 587014 581703 587016
rect 581637 587011 581703 587014
rect -960 580002 480 580092
rect 2037 580002 2103 580005
rect -960 580000 2103 580002
rect -960 579944 2042 580000
rect 2098 579944 2103 580000
rect -960 579942 2103 579944
rect -960 579852 480 579942
rect 2037 579939 2103 579942
rect 581637 577690 581703 577693
rect 583520 577690 584960 577780
rect 581637 577688 584960 577690
rect 581637 577632 581642 577688
rect 581698 577632 584960 577688
rect 581637 577630 584960 577632
rect 581637 577627 581703 577630
rect 583520 577540 584960 577630
rect 2037 575786 2103 575789
rect 2037 575784 3220 575786
rect 2037 575728 2042 575784
rect 2098 575728 3220 575784
rect 2037 575726 3220 575728
rect 2037 575723 2103 575726
rect 581637 574018 581703 574021
rect 580796 574016 581703 574018
rect 580796 573960 581642 574016
rect 581698 573960 581703 574016
rect 580796 573958 581703 573960
rect 581637 573955 581703 573958
rect -960 566946 480 567036
rect 1485 566946 1551 566949
rect -960 566944 1551 566946
rect -960 566888 1490 566944
rect 1546 566888 1551 566944
rect -960 566886 1551 566888
rect -960 566796 480 566886
rect 1485 566883 1551 566886
rect 582373 564362 582439 564365
rect 583520 564362 584960 564452
rect 582373 564360 584960 564362
rect 582373 564304 582378 564360
rect 582434 564304 584960 564360
rect 582373 564302 584960 564304
rect 582373 564299 582439 564302
rect 583520 564212 584960 564302
rect 1485 563002 1551 563005
rect 1485 563000 3220 563002
rect 1485 562944 1490 563000
rect 1546 562944 3220 563000
rect 1485 562942 3220 562944
rect 1485 562939 1551 562942
rect 582373 560962 582439 560965
rect 580796 560960 582439 560962
rect 580796 560904 582378 560960
rect 582434 560904 582439 560960
rect 580796 560902 582439 560904
rect 582373 560899 582439 560902
rect -960 553890 480 553980
rect 1485 553890 1551 553893
rect -960 553888 1551 553890
rect -960 553832 1490 553888
rect 1546 553832 1551 553888
rect -960 553830 1551 553832
rect -960 553740 480 553830
rect 1485 553827 1551 553830
rect 581637 551170 581703 551173
rect 583520 551170 584960 551260
rect 581637 551168 584960 551170
rect 581637 551112 581642 551168
rect 581698 551112 584960 551168
rect 581637 551110 584960 551112
rect 581637 551107 581703 551110
rect 583520 551020 584960 551110
rect 1485 550218 1551 550221
rect 1485 550216 3220 550218
rect 1485 550160 1490 550216
rect 1546 550160 3220 550216
rect 1485 550158 3220 550160
rect 1485 550155 1551 550158
rect 581637 547770 581703 547773
rect 580796 547768 581703 547770
rect 580796 547712 581642 547768
rect 581698 547712 581703 547768
rect 580796 547710 581703 547712
rect 581637 547707 581703 547710
rect -960 540834 480 540924
rect 1393 540834 1459 540837
rect -960 540832 1459 540834
rect -960 540776 1398 540832
rect 1454 540776 1459 540832
rect -960 540774 1459 540776
rect -960 540684 480 540774
rect 1393 540771 1459 540774
rect 582373 537842 582439 537845
rect 583520 537842 584960 537932
rect 582373 537840 584960 537842
rect 582373 537784 582378 537840
rect 582434 537784 584960 537840
rect 582373 537782 584960 537784
rect 582373 537779 582439 537782
rect 583520 537692 584960 537782
rect 1393 537434 1459 537437
rect 1393 537432 3220 537434
rect 1393 537376 1398 537432
rect 1454 537376 3220 537432
rect 1393 537374 3220 537376
rect 1393 537371 1459 537374
rect 582373 534850 582439 534853
rect 580796 534848 582439 534850
rect 580796 534792 582378 534848
rect 582434 534792 582439 534848
rect 580796 534790 582439 534792
rect 582373 534787 582439 534790
rect -960 527914 480 528004
rect 1485 527914 1551 527917
rect -960 527912 1551 527914
rect -960 527856 1490 527912
rect 1546 527856 1551 527912
rect -960 527854 1551 527856
rect -960 527764 480 527854
rect 1485 527851 1551 527854
rect 1485 524650 1551 524653
rect 1485 524648 3220 524650
rect 1485 524592 1490 524648
rect 1546 524592 3220 524648
rect 1485 524590 3220 524592
rect 1485 524587 1551 524590
rect 582373 524514 582439 524517
rect 583520 524514 584960 524604
rect 582373 524512 584960 524514
rect 582373 524456 582378 524512
rect 582434 524456 584960 524512
rect 582373 524454 584960 524456
rect 582373 524451 582439 524454
rect 583520 524364 584960 524454
rect 582373 521794 582439 521797
rect 580796 521792 582439 521794
rect 580796 521736 582378 521792
rect 582434 521736 582439 521792
rect 580796 521734 582439 521736
rect 582373 521731 582439 521734
rect -960 514858 480 514948
rect 1577 514858 1643 514861
rect -960 514856 1643 514858
rect -960 514800 1582 514856
rect 1638 514800 1643 514856
rect -960 514798 1643 514800
rect -960 514708 480 514798
rect 1577 514795 1643 514798
rect 1577 511866 1643 511869
rect 1577 511864 3220 511866
rect 1577 511808 1582 511864
rect 1638 511808 3220 511864
rect 1577 511806 3220 511808
rect 1577 511803 1643 511806
rect 582373 511322 582439 511325
rect 583520 511322 584960 511412
rect 582373 511320 584960 511322
rect 582373 511264 582378 511320
rect 582434 511264 584960 511320
rect 582373 511262 584960 511264
rect 582373 511259 582439 511262
rect 583520 511172 584960 511262
rect 582373 508738 582439 508741
rect 580796 508736 582439 508738
rect 580796 508680 582378 508736
rect 582434 508680 582439 508736
rect 580796 508678 582439 508680
rect 582373 508675 582439 508678
rect -960 501802 480 501892
rect 1577 501802 1643 501805
rect -960 501800 1643 501802
rect -960 501744 1582 501800
rect 1638 501744 1643 501800
rect -960 501742 1643 501744
rect -960 501652 480 501742
rect 1577 501739 1643 501742
rect 1577 499082 1643 499085
rect 1577 499080 3220 499082
rect 1577 499024 1582 499080
rect 1638 499024 3220 499080
rect 1577 499022 3220 499024
rect 1577 499019 1643 499022
rect 581637 497994 581703 497997
rect 583520 497994 584960 498084
rect 581637 497992 584960 497994
rect 581637 497936 581642 497992
rect 581698 497936 584960 497992
rect 581637 497934 584960 497936
rect 581637 497931 581703 497934
rect 583520 497844 584960 497934
rect 581637 495682 581703 495685
rect 580796 495680 581703 495682
rect 580796 495624 581642 495680
rect 581698 495624 581703 495680
rect 580796 495622 581703 495624
rect 581637 495619 581703 495622
rect -960 488746 480 488836
rect 1577 488746 1643 488749
rect -960 488744 1643 488746
rect -960 488688 1582 488744
rect 1638 488688 1643 488744
rect -960 488686 1643 488688
rect -960 488596 480 488686
rect 1577 488683 1643 488686
rect 1577 486298 1643 486301
rect 1577 486296 3220 486298
rect 1577 486240 1582 486296
rect 1638 486240 3220 486296
rect 1577 486238 3220 486240
rect 1577 486235 1643 486238
rect 582373 484666 582439 484669
rect 583520 484666 584960 484756
rect 582373 484664 584960 484666
rect 582373 484608 582378 484664
rect 582434 484608 584960 484664
rect 582373 484606 584960 484608
rect 582373 484603 582439 484606
rect 583520 484516 584960 484606
rect 582373 482626 582439 482629
rect 580796 482624 582439 482626
rect 580796 482568 582378 482624
rect 582434 482568 582439 482624
rect 580796 482566 582439 482568
rect 582373 482563 582439 482566
rect -960 475690 480 475780
rect 2773 475690 2839 475693
rect -960 475688 2839 475690
rect -960 475632 2778 475688
rect 2834 475632 2839 475688
rect -960 475630 2839 475632
rect -960 475540 480 475630
rect 2773 475627 2839 475630
rect 2773 473514 2839 473517
rect 2773 473512 3220 473514
rect 2773 473456 2778 473512
rect 2834 473456 3220 473512
rect 2773 473454 3220 473456
rect 2773 473451 2839 473454
rect 581637 471474 581703 471477
rect 583520 471474 584960 471564
rect 581637 471472 584960 471474
rect 581637 471416 581642 471472
rect 581698 471416 584960 471472
rect 581637 471414 584960 471416
rect 581637 471411 581703 471414
rect 583520 471324 584960 471414
rect 581637 469570 581703 469573
rect 580796 469568 581703 469570
rect 580796 469512 581642 469568
rect 581698 469512 581703 469568
rect 580796 469510 581703 469512
rect 581637 469507 581703 469510
rect -960 462634 480 462724
rect 1577 462634 1643 462637
rect -960 462632 1643 462634
rect -960 462576 1582 462632
rect 1638 462576 1643 462632
rect -960 462574 1643 462576
rect -960 462484 480 462574
rect 1577 462571 1643 462574
rect 1577 460730 1643 460733
rect 1577 460728 3220 460730
rect 1577 460672 1582 460728
rect 1638 460672 3220 460728
rect 1577 460670 3220 460672
rect 1577 460667 1643 460670
rect 581637 458146 581703 458149
rect 583520 458146 584960 458236
rect 581637 458144 584960 458146
rect 581637 458088 581642 458144
rect 581698 458088 584960 458144
rect 581637 458086 584960 458088
rect 581637 458083 581703 458086
rect 583520 457996 584960 458086
rect 581637 456514 581703 456517
rect 580796 456512 581703 456514
rect 580796 456456 581642 456512
rect 581698 456456 581703 456512
rect 580796 456454 581703 456456
rect 581637 456451 581703 456454
rect -960 449578 480 449668
rect 2773 449578 2839 449581
rect -960 449576 2839 449578
rect -960 449520 2778 449576
rect 2834 449520 2839 449576
rect -960 449518 2839 449520
rect -960 449428 480 449518
rect 2773 449515 2839 449518
rect 2773 447946 2839 447949
rect 2773 447944 3220 447946
rect 2773 447888 2778 447944
rect 2834 447888 3220 447944
rect 2773 447886 3220 447888
rect 2773 447883 2839 447886
rect 583520 444818 584960 444908
rect 583342 444758 584960 444818
rect 583342 444682 583402 444758
rect 583520 444682 584960 444758
rect 583342 444668 584960 444682
rect 583342 444622 583586 444668
rect 583526 444138 583586 444622
rect 580766 444078 583586 444138
rect 580766 443428 580826 444078
rect -960 436658 480 436748
rect 2773 436658 2839 436661
rect -960 436656 2839 436658
rect -960 436600 2778 436656
rect 2834 436600 2839 436656
rect -960 436598 2839 436600
rect -960 436508 480 436598
rect 2773 436595 2839 436598
rect 2773 435162 2839 435165
rect 2773 435160 3220 435162
rect 2773 435104 2778 435160
rect 2834 435104 3220 435160
rect 2773 435102 3220 435104
rect 2773 435099 2839 435102
rect 583520 431626 584960 431716
rect 583342 431566 584960 431626
rect 583342 431490 583402 431566
rect 583520 431490 584960 431566
rect 583342 431476 584960 431490
rect 583342 431430 583586 431476
rect 583526 431082 583586 431430
rect 580766 431022 583586 431082
rect 580766 430372 580826 431022
rect -960 423602 480 423692
rect 2773 423602 2839 423605
rect -960 423600 2839 423602
rect -960 423544 2778 423600
rect 2834 423544 2839 423600
rect -960 423542 2839 423544
rect -960 423452 480 423542
rect 2773 423539 2839 423542
rect 2773 422378 2839 422381
rect 2773 422376 3220 422378
rect 2773 422320 2778 422376
rect 2834 422320 3220 422376
rect 2773 422318 3220 422320
rect 2773 422315 2839 422318
rect 583520 418298 584960 418388
rect 583342 418238 584960 418298
rect 583342 418162 583402 418238
rect 583520 418162 584960 418238
rect 583342 418148 584960 418162
rect 583342 418102 583586 418148
rect 583526 417754 583586 418102
rect 580766 417694 583586 417754
rect 580766 417316 580826 417694
rect -960 410546 480 410636
rect -960 410486 3250 410546
rect -960 410396 480 410486
rect 3190 409564 3250 410486
rect 583520 404970 584960 405060
rect 580766 404910 584960 404970
rect 580766 404260 580826 404910
rect 583520 404820 584960 404910
rect -960 397490 480 397580
rect -960 397430 3250 397490
rect -960 397340 480 397430
rect 3190 396780 3250 397430
rect 583520 391778 584960 391868
rect 580766 391718 584960 391778
rect 580766 391204 580826 391718
rect 583520 391628 584960 391718
rect -960 384434 480 384524
rect -960 384374 3250 384434
rect -960 384284 480 384374
rect 3190 383996 3250 384374
rect 583520 378450 584960 378540
rect 580766 378390 584960 378450
rect 580766 378148 580826 378390
rect 583520 378300 584960 378390
rect -960 371378 480 371468
rect -960 371318 3250 371378
rect -960 371228 480 371318
rect 3190 371212 3250 371318
rect 583520 365122 584960 365212
rect 580796 365062 584960 365122
rect 583520 364972 584960 365062
rect -960 358458 480 358548
rect -960 358398 3220 358458
rect -960 358308 480 358398
rect 583520 351930 584960 352020
rect 580796 351870 584960 351930
rect 583520 351780 584960 351870
rect -960 345402 480 345492
rect 1534 345478 3220 345538
rect 1534 345402 1594 345478
rect -960 345342 1594 345402
rect -960 345252 480 345342
rect 580766 338602 580826 338844
rect 583520 338602 584960 338692
rect 580766 338542 584960 338602
rect 583520 338452 584960 338542
rect -960 332346 480 332436
rect 3190 332346 3250 332724
rect -960 332286 3250 332346
rect -960 332196 480 332286
rect 580766 325274 580826 325788
rect 583520 325274 584960 325364
rect 580766 325214 584960 325274
rect 583520 325124 584960 325214
rect -960 319290 480 319380
rect 3190 319290 3250 319940
rect -960 319230 3250 319290
rect -960 319140 480 319230
rect 580766 312082 580826 312732
rect 583520 312082 584960 312172
rect 580766 312022 584960 312082
rect 583520 311932 584960 312022
rect -960 306234 480 306324
rect 3190 306234 3250 307156
rect -960 306174 3250 306234
rect -960 306084 480 306174
rect 580766 299298 580826 299676
rect 580766 299238 583586 299298
rect 583526 298890 583586 299238
rect 583342 298844 583586 298890
rect 583342 298830 584960 298844
rect 583342 298754 583402 298830
rect 583520 298754 584960 298830
rect 583342 298694 584960 298754
rect 583520 298604 584960 298694
rect 1301 294402 1367 294405
rect 1301 294400 3220 294402
rect 1301 294344 1306 294400
rect 1362 294344 3220 294400
rect 1301 294342 3220 294344
rect 1301 294339 1367 294342
rect -960 293178 480 293268
rect 1301 293178 1367 293181
rect -960 293176 1367 293178
rect -960 293120 1306 293176
rect 1362 293120 1367 293176
rect -960 293118 1367 293120
rect -960 293028 480 293118
rect 1301 293115 1367 293118
rect 580766 285970 580826 286620
rect 580766 285910 583586 285970
rect 583526 285562 583586 285910
rect 583342 285516 583586 285562
rect 583342 285502 584960 285516
rect 583342 285426 583402 285502
rect 583520 285426 584960 285502
rect 583342 285366 584960 285426
rect 583520 285276 584960 285366
rect 2773 281618 2839 281621
rect 2773 281616 3220 281618
rect 2773 281560 2778 281616
rect 2834 281560 3220 281616
rect 2773 281558 3220 281560
rect 2773 281555 2839 281558
rect -960 280122 480 280212
rect 2773 280122 2839 280125
rect -960 280120 2839 280122
rect -960 280064 2778 280120
rect 2834 280064 2839 280120
rect -960 280062 2839 280064
rect -960 279972 480 280062
rect 2773 280059 2839 280062
rect 580766 272914 580826 273564
rect 580766 272854 583586 272914
rect 583526 272370 583586 272854
rect 583342 272324 583586 272370
rect 583342 272310 584960 272324
rect 583342 272234 583402 272310
rect 583520 272234 584960 272310
rect 583342 272174 584960 272234
rect 583520 272084 584960 272174
rect 1301 268834 1367 268837
rect 1301 268832 3220 268834
rect 1301 268776 1306 268832
rect 1362 268776 3220 268832
rect 1301 268774 3220 268776
rect 1301 268771 1367 268774
rect -960 267202 480 267292
rect 1301 267202 1367 267205
rect -960 267200 1367 267202
rect -960 267144 1306 267200
rect 1362 267144 1367 267200
rect -960 267142 1367 267144
rect -960 267052 480 267142
rect 1301 267139 1367 267142
rect 582373 260538 582439 260541
rect 580796 260536 582439 260538
rect 580796 260480 582378 260536
rect 582434 260480 582439 260536
rect 580796 260478 582439 260480
rect 582373 260475 582439 260478
rect 582373 258906 582439 258909
rect 583520 258906 584960 258996
rect 582373 258904 584960 258906
rect 582373 258848 582378 258904
rect 582434 258848 584960 258904
rect 582373 258846 584960 258848
rect 582373 258843 582439 258846
rect 583520 258756 584960 258846
rect 1301 256050 1367 256053
rect 1301 256048 3220 256050
rect 1301 255992 1306 256048
rect 1362 255992 3220 256048
rect 1301 255990 3220 255992
rect 1301 255987 1367 255990
rect -960 254146 480 254236
rect 1301 254146 1367 254149
rect -960 254144 1367 254146
rect -960 254088 1306 254144
rect 1362 254088 1367 254144
rect -960 254086 1367 254088
rect -960 253996 480 254086
rect 1301 254083 1367 254086
rect 580766 247074 580826 247452
rect 580901 247074 580967 247077
rect 580766 247072 580967 247074
rect 580766 247016 580906 247072
rect 580962 247016 580967 247072
rect 580766 247014 580967 247016
rect 580901 247011 580967 247014
rect 580901 245578 580967 245581
rect 583520 245578 584960 245668
rect 580901 245576 584960 245578
rect 580901 245520 580906 245576
rect 580962 245520 584960 245576
rect 580901 245518 584960 245520
rect 580901 245515 580967 245518
rect 583520 245428 584960 245518
rect 2773 243266 2839 243269
rect 2773 243264 3220 243266
rect 2773 243208 2778 243264
rect 2834 243208 3220 243264
rect 2773 243206 3220 243208
rect 2773 243203 2839 243206
rect -960 241090 480 241180
rect 2773 241090 2839 241093
rect -960 241088 2839 241090
rect -960 241032 2778 241088
rect 2834 241032 2839 241088
rect -960 241030 2839 241032
rect -960 240940 480 241030
rect 2773 241027 2839 241030
rect 582373 234426 582439 234429
rect 580796 234424 582439 234426
rect 580796 234368 582378 234424
rect 582434 234368 582439 234424
rect 580796 234366 582439 234368
rect 582373 234363 582439 234366
rect 582373 232386 582439 232389
rect 583520 232386 584960 232476
rect 582373 232384 584960 232386
rect 582373 232328 582378 232384
rect 582434 232328 584960 232384
rect 582373 232326 584960 232328
rect 582373 232323 582439 232326
rect 583520 232236 584960 232326
rect 2773 230618 2839 230621
rect 2773 230616 3220 230618
rect 2773 230560 2778 230616
rect 2834 230560 3220 230616
rect 2773 230558 3220 230560
rect 2773 230555 2839 230558
rect -960 228034 480 228124
rect 2773 228034 2839 228037
rect -960 228032 2839 228034
rect -960 227976 2778 228032
rect 2834 227976 2839 228032
rect -960 227974 2839 227976
rect -960 227884 480 227974
rect 2773 227971 2839 227974
rect 580766 220962 580826 221340
rect 580901 220962 580967 220965
rect 580766 220960 580967 220962
rect 580766 220904 580906 220960
rect 580962 220904 580967 220960
rect 580766 220902 580967 220904
rect 580901 220899 580967 220902
rect 580901 219058 580967 219061
rect 583520 219058 584960 219148
rect 580901 219056 584960 219058
rect 580901 219000 580906 219056
rect 580962 219000 584960 219056
rect 580901 218998 584960 219000
rect 580901 218995 580967 218998
rect 583520 218908 584960 218998
rect 2773 217698 2839 217701
rect 2773 217696 3220 217698
rect 2773 217640 2778 217696
rect 2834 217640 3220 217696
rect 2773 217638 3220 217640
rect 2773 217635 2839 217638
rect -960 214978 480 215068
rect 2773 214978 2839 214981
rect -960 214976 2839 214978
rect -960 214920 2778 214976
rect 2834 214920 2839 214976
rect -960 214918 2839 214920
rect -960 214828 480 214918
rect 2773 214915 2839 214918
rect 582373 208314 582439 208317
rect 580796 208312 582439 208314
rect 580796 208256 582378 208312
rect 582434 208256 582439 208312
rect 580796 208254 582439 208256
rect 582373 208251 582439 208254
rect 582373 205730 582439 205733
rect 583520 205730 584960 205820
rect 582373 205728 584960 205730
rect 582373 205672 582378 205728
rect 582434 205672 584960 205728
rect 582373 205670 584960 205672
rect 582373 205667 582439 205670
rect 583520 205580 584960 205670
rect 2773 204914 2839 204917
rect 2773 204912 3220 204914
rect 2773 204856 2778 204912
rect 2834 204856 3220 204912
rect 2773 204854 3220 204856
rect 2773 204851 2839 204854
rect -960 201922 480 202012
rect 2773 201922 2839 201925
rect -960 201920 2839 201922
rect -960 201864 2778 201920
rect 2834 201864 2839 201920
rect -960 201862 2839 201864
rect -960 201772 480 201862
rect 2773 201859 2839 201862
rect 580766 194714 580826 195228
rect 580901 194714 580967 194717
rect 580766 194712 580967 194714
rect 580766 194656 580906 194712
rect 580962 194656 580967 194712
rect 580766 194654 580967 194656
rect 580901 194651 580967 194654
rect 580901 192538 580967 192541
rect 583520 192538 584960 192628
rect 580901 192536 584960 192538
rect 580901 192480 580906 192536
rect 580962 192480 584960 192536
rect 580901 192478 584960 192480
rect 580901 192475 580967 192478
rect 583520 192388 584960 192478
rect 1301 192130 1367 192133
rect 1301 192128 3220 192130
rect 1301 192072 1306 192128
rect 1362 192072 3220 192128
rect 1301 192070 3220 192072
rect 1301 192067 1367 192070
rect -960 188866 480 188956
rect 1301 188866 1367 188869
rect -960 188864 1367 188866
rect -960 188808 1306 188864
rect 1362 188808 1367 188864
rect -960 188806 1367 188808
rect -960 188716 480 188806
rect 1301 188803 1367 188806
rect 580901 182474 580967 182477
rect 580766 182472 580967 182474
rect 580766 182416 580906 182472
rect 580962 182416 580967 182472
rect 580766 182414 580967 182416
rect 580766 182308 580826 182414
rect 580901 182411 580967 182414
rect 2773 179346 2839 179349
rect 2773 179344 3220 179346
rect 2773 179288 2778 179344
rect 2834 179288 3220 179344
rect 2773 179286 3220 179288
rect 2773 179283 2839 179286
rect 580901 179210 580967 179213
rect 583520 179210 584960 179300
rect 580901 179208 584960 179210
rect 580901 179152 580906 179208
rect 580962 179152 584960 179208
rect 580901 179150 584960 179152
rect 580901 179147 580967 179150
rect 583520 179060 584960 179150
rect -960 175946 480 176036
rect 2773 175946 2839 175949
rect -960 175944 2839 175946
rect -960 175888 2778 175944
rect 2834 175888 2839 175944
rect -960 175886 2839 175888
rect -960 175796 480 175886
rect 2773 175883 2839 175886
rect 580766 168602 580826 169116
rect 580901 168602 580967 168605
rect 580766 168600 580967 168602
rect 580766 168544 580906 168600
rect 580962 168544 580967 168600
rect 580766 168542 580967 168544
rect 580901 168539 580967 168542
rect 2773 166562 2839 166565
rect 2773 166560 3220 166562
rect 2773 166504 2778 166560
rect 2834 166504 3220 166560
rect 2773 166502 3220 166504
rect 2773 166499 2839 166502
rect 580901 165882 580967 165885
rect 583520 165882 584960 165972
rect 580901 165880 584960 165882
rect 580901 165824 580906 165880
rect 580962 165824 584960 165880
rect 580901 165822 584960 165824
rect 580901 165819 580967 165822
rect 583520 165732 584960 165822
rect -960 162890 480 162980
rect 2773 162890 2839 162893
rect -960 162888 2839 162890
rect -960 162832 2778 162888
rect 2834 162832 2839 162888
rect -960 162830 2839 162832
rect -960 162740 480 162830
rect 2773 162827 2839 162830
rect 580901 156362 580967 156365
rect 580766 156360 580967 156362
rect 580766 156304 580906 156360
rect 580962 156304 580967 156360
rect 580766 156302 580967 156304
rect 580766 156196 580826 156302
rect 580901 156299 580967 156302
rect 1301 153778 1367 153781
rect 1301 153776 3220 153778
rect 1301 153720 1306 153776
rect 1362 153720 3220 153776
rect 1301 153718 3220 153720
rect 1301 153715 1367 153718
rect 580901 152690 580967 152693
rect 583520 152690 584960 152780
rect 580901 152688 584960 152690
rect 580901 152632 580906 152688
rect 580962 152632 584960 152688
rect 580901 152630 584960 152632
rect 580901 152627 580967 152630
rect 583520 152540 584960 152630
rect -960 149834 480 149924
rect 1301 149834 1367 149837
rect -960 149832 1367 149834
rect -960 149776 1306 149832
rect 1362 149776 1367 149832
rect -960 149774 1367 149776
rect -960 149684 480 149774
rect 1301 149771 1367 149774
rect 580766 142626 580826 143004
rect 580901 142626 580967 142629
rect 580766 142624 580967 142626
rect 580766 142568 580906 142624
rect 580962 142568 580967 142624
rect 580766 142566 580967 142568
rect 580901 142563 580967 142566
rect 565 140994 631 140997
rect 565 140992 3220 140994
rect 565 140936 570 140992
rect 626 140936 3220 140992
rect 565 140934 3220 140936
rect 565 140931 631 140934
rect 580901 139362 580967 139365
rect 583520 139362 584960 139452
rect 580901 139360 584960 139362
rect 580901 139304 580906 139360
rect 580962 139304 584960 139360
rect 580901 139302 584960 139304
rect 580901 139299 580967 139302
rect 583520 139212 584960 139302
rect -960 136778 480 136868
rect 565 136778 631 136781
rect -960 136776 631 136778
rect -960 136720 570 136776
rect 626 136720 631 136776
rect -960 136718 631 136720
rect -960 136628 480 136718
rect 565 136715 631 136718
rect 580901 130250 580967 130253
rect 580766 130248 580967 130250
rect 580766 130192 580906 130248
rect 580962 130192 580967 130248
rect 580766 130190 580967 130192
rect 580766 130084 580826 130190
rect 580901 130187 580967 130190
rect 749 128210 815 128213
rect 749 128208 3220 128210
rect 749 128152 754 128208
rect 810 128152 3220 128208
rect 749 128150 3220 128152
rect 749 128147 815 128150
rect 580901 126034 580967 126037
rect 583520 126034 584960 126124
rect 580901 126032 584960 126034
rect 580901 125976 580906 126032
rect 580962 125976 584960 126032
rect 580901 125974 584960 125976
rect 580901 125971 580967 125974
rect 583520 125884 584960 125974
rect -960 123722 480 123812
rect 749 123722 815 123725
rect -960 123720 815 123722
rect -960 123664 754 123720
rect 810 123664 815 123720
rect -960 123662 815 123664
rect -960 123572 480 123662
rect 749 123659 815 123662
rect 579889 116378 579955 116381
rect 580030 116378 580090 116892
rect 579889 116376 580090 116378
rect 579889 116320 579894 116376
rect 579950 116320 580090 116376
rect 579889 116318 580090 116320
rect 579889 116315 579955 116318
rect 1301 115426 1367 115429
rect 1301 115424 3220 115426
rect 1301 115368 1306 115424
rect 1362 115368 3220 115424
rect 1301 115366 3220 115368
rect 1301 115363 1367 115366
rect 579889 112842 579955 112845
rect 583520 112842 584960 112932
rect 579889 112840 584960 112842
rect 579889 112784 579894 112840
rect 579950 112784 584960 112840
rect 579889 112782 584960 112784
rect 579889 112779 579955 112782
rect 583520 112692 584960 112782
rect -960 110666 480 110756
rect 1301 110666 1367 110669
rect -960 110664 1367 110666
rect -960 110608 1306 110664
rect 1362 110608 1367 110664
rect -960 110606 1367 110608
rect -960 110516 480 110606
rect 1301 110603 1367 110606
rect 580766 103594 580826 103836
rect 580901 103594 580967 103597
rect 580766 103592 580967 103594
rect 580766 103536 580906 103592
rect 580962 103536 580967 103592
rect 580766 103534 580967 103536
rect 580901 103531 580967 103534
rect 1577 102642 1643 102645
rect 1577 102640 3220 102642
rect 1577 102584 1582 102640
rect 1638 102584 3220 102640
rect 1577 102582 3220 102584
rect 1577 102579 1643 102582
rect 580901 99514 580967 99517
rect 583520 99514 584960 99604
rect 580901 99512 584960 99514
rect 580901 99456 580906 99512
rect 580962 99456 584960 99512
rect 580901 99454 584960 99456
rect 580901 99451 580967 99454
rect 583520 99364 584960 99454
rect -960 97610 480 97700
rect 1577 97610 1643 97613
rect -960 97608 1643 97610
rect -960 97552 1582 97608
rect 1638 97552 1643 97608
rect -960 97550 1643 97552
rect -960 97460 480 97550
rect 1577 97547 1643 97550
rect 580766 90266 580826 90780
rect 580901 90266 580967 90269
rect 580766 90264 580967 90266
rect 580766 90208 580906 90264
rect 580962 90208 580967 90264
rect 580766 90206 580967 90208
rect 580901 90203 580967 90206
rect 1577 89858 1643 89861
rect 1577 89856 3220 89858
rect 1577 89800 1582 89856
rect 1638 89800 3220 89856
rect 1577 89798 3220 89800
rect 1577 89795 1643 89798
rect 580901 86186 580967 86189
rect 583520 86186 584960 86276
rect 580901 86184 584960 86186
rect 580901 86128 580906 86184
rect 580962 86128 584960 86184
rect 580901 86126 584960 86128
rect 580901 86123 580967 86126
rect 583520 86036 584960 86126
rect -960 84690 480 84780
rect 1577 84690 1643 84693
rect -960 84688 1643 84690
rect -960 84632 1582 84688
rect 1638 84632 1643 84688
rect -960 84630 1643 84632
rect -960 84540 480 84630
rect 1577 84627 1643 84630
rect 579889 77346 579955 77349
rect 580030 77346 580090 77724
rect 579889 77344 580090 77346
rect 579889 77288 579894 77344
rect 579950 77288 580090 77344
rect 579889 77286 580090 77288
rect 579889 77283 579955 77286
rect 1577 77074 1643 77077
rect 1577 77072 3220 77074
rect 1577 77016 1582 77072
rect 1638 77016 3220 77072
rect 1577 77014 3220 77016
rect 1577 77011 1643 77014
rect 579889 72994 579955 72997
rect 583520 72994 584960 73084
rect 579889 72992 584960 72994
rect 579889 72936 579894 72992
rect 579950 72936 584960 72992
rect 579889 72934 584960 72936
rect 579889 72931 579955 72934
rect 583520 72844 584960 72934
rect -960 71634 480 71724
rect 1577 71634 1643 71637
rect -960 71632 1643 71634
rect -960 71576 1582 71632
rect 1638 71576 1643 71632
rect -960 71574 1643 71576
rect -960 71484 480 71574
rect 1577 71571 1643 71574
rect 1485 64290 1551 64293
rect 1485 64288 3220 64290
rect 1485 64232 1490 64288
rect 1546 64232 3220 64288
rect 1485 64230 3220 64232
rect 1485 64227 1551 64230
rect 580766 64154 580826 64668
rect 580901 64154 580967 64157
rect 580766 64152 580967 64154
rect 580766 64096 580906 64152
rect 580962 64096 580967 64152
rect 580766 64094 580967 64096
rect 580901 64091 580967 64094
rect 580901 59666 580967 59669
rect 583520 59666 584960 59756
rect 580901 59664 584960 59666
rect 580901 59608 580906 59664
rect 580962 59608 584960 59664
rect 580901 59606 584960 59608
rect 580901 59603 580967 59606
rect 583520 59516 584960 59606
rect -960 58578 480 58668
rect 1485 58578 1551 58581
rect -960 58576 1551 58578
rect -960 58520 1490 58576
rect 1546 58520 1551 58576
rect -960 58518 1551 58520
rect -960 58428 480 58518
rect 1485 58515 1551 58518
rect 2037 51506 2103 51509
rect 2037 51504 3220 51506
rect 2037 51448 2042 51504
rect 2098 51448 3220 51504
rect 2037 51446 3220 51448
rect 2037 51443 2103 51446
rect 580766 51098 580826 51612
rect 580901 51098 580967 51101
rect 580766 51096 580967 51098
rect 580766 51040 580906 51096
rect 580962 51040 580967 51096
rect 580766 51038 580967 51040
rect 580901 51035 580967 51038
rect 580901 46338 580967 46341
rect 583520 46338 584960 46428
rect 580901 46336 584960 46338
rect 580901 46280 580906 46336
rect 580962 46280 584960 46336
rect 580901 46278 584960 46280
rect 580901 46275 580967 46278
rect 583520 46188 584960 46278
rect -960 45522 480 45612
rect 2037 45522 2103 45525
rect -960 45520 2103 45522
rect -960 45464 2042 45520
rect 2098 45464 2103 45520
rect -960 45462 2103 45464
rect -960 45372 480 45462
rect 2037 45459 2103 45462
rect 2037 38722 2103 38725
rect 2037 38720 3220 38722
rect 2037 38664 2042 38720
rect 2098 38664 3220 38720
rect 2037 38662 3220 38664
rect 2037 38659 2103 38662
rect 580766 38042 580826 38556
rect 580901 38042 580967 38045
rect 580766 38040 580967 38042
rect 580766 37984 580906 38040
rect 580962 37984 580967 38040
rect 580766 37982 580967 37984
rect 580901 37979 580967 37982
rect 580901 33146 580967 33149
rect 583520 33146 584960 33236
rect 580901 33144 584960 33146
rect 580901 33088 580906 33144
rect 580962 33088 584960 33144
rect 580901 33086 584960 33088
rect 580901 33083 580967 33086
rect 583520 32996 584960 33086
rect -960 32466 480 32556
rect 2037 32466 2103 32469
rect -960 32464 2103 32466
rect -960 32408 2042 32464
rect 2098 32408 2103 32464
rect -960 32406 2103 32408
rect -960 32316 480 32406
rect 2037 32403 2103 32406
rect 1485 25938 1551 25941
rect 1485 25936 3220 25938
rect 1485 25880 1490 25936
rect 1546 25880 3220 25936
rect 1485 25878 3220 25880
rect 1485 25875 1551 25878
rect 580766 24986 580826 25500
rect 580901 24986 580967 24989
rect 580766 24984 580967 24986
rect 580766 24928 580906 24984
rect 580962 24928 580967 24984
rect 580766 24926 580967 24928
rect 580901 24923 580967 24926
rect 580901 19818 580967 19821
rect 583520 19818 584960 19908
rect 580901 19816 584960 19818
rect 580901 19760 580906 19816
rect 580962 19760 584960 19816
rect 580901 19758 584960 19760
rect 580901 19755 580967 19758
rect 583520 19668 584960 19758
rect -960 19410 480 19500
rect 1485 19410 1551 19413
rect -960 19408 1551 19410
rect -960 19352 1490 19408
rect 1546 19352 1551 19408
rect -960 19350 1551 19352
rect -960 19260 480 19350
rect 1485 19347 1551 19350
rect 2037 13154 2103 13157
rect 2037 13152 3220 13154
rect 2037 13096 2042 13152
rect 2098 13096 3220 13152
rect 2037 13094 3220 13096
rect 2037 13091 2103 13094
rect 582373 12474 582439 12477
rect 580796 12472 582439 12474
rect 580796 12416 582378 12472
rect 582434 12416 582439 12472
rect 580796 12414 582439 12416
rect 582373 12411 582439 12414
rect 582373 6626 582439 6629
rect 583520 6626 584960 6716
rect 582373 6624 584960 6626
rect -960 6490 480 6580
rect 582373 6568 582378 6624
rect 582434 6568 584960 6624
rect 582373 6566 584960 6568
rect 582373 6563 582439 6566
rect 2037 6490 2103 6493
rect -960 6488 2103 6490
rect -960 6432 2042 6488
rect 2098 6432 2103 6488
rect 583520 6476 584960 6566
rect -960 6430 2103 6432
rect -960 6340 480 6430
rect 2037 6427 2103 6430
rect 28901 642 28967 645
rect 46289 642 46355 645
rect 28901 640 46355 642
rect 28901 584 28906 640
rect 28962 584 46294 640
rect 46350 584 46355 640
rect 28901 582 46355 584
rect 28901 579 28967 582
rect 46289 579 46355 582
rect 12157 506 12223 509
rect 30833 506 30899 509
rect 12157 504 30899 506
rect 12157 448 12162 504
rect 12218 448 30838 504
rect 30894 448 30899 504
rect 12157 446 30899 448
rect 12157 443 12223 446
rect 30833 443 30899 446
rect 13721 370 13787 373
rect 31937 370 32003 373
rect 13721 368 32003 370
rect 13721 312 13726 368
rect 13782 312 31942 368
rect 31998 312 32003 368
rect 13721 310 32003 312
rect 13721 307 13787 310
rect 31937 307 32003 310
rect 6269 234 6335 237
rect 25037 234 25103 237
rect 6269 232 25103 234
rect 6269 176 6274 232
rect 6330 176 25042 232
rect 25098 176 25103 232
rect 6269 174 25103 176
rect 6269 171 6335 174
rect 25037 171 25103 174
rect 25681 234 25747 237
rect 42701 234 42767 237
rect 25681 232 42767 234
rect 25681 176 25686 232
rect 25742 176 42706 232
rect 42762 176 42767 232
rect 25681 174 42767 176
rect 25681 171 25747 174
rect 42701 171 42767 174
rect 46841 234 46907 237
rect 62849 234 62915 237
rect 46841 232 62915 234
rect 46841 176 46846 232
rect 46902 176 62854 232
rect 62910 176 62915 232
rect 46841 174 62915 176
rect 46841 171 46907 174
rect 62849 171 62915 174
rect 5441 98 5507 101
rect 23933 98 23999 101
rect 5441 96 23999 98
rect 5441 40 5446 96
rect 5502 40 23938 96
rect 23994 40 23999 96
rect 5441 38 23999 40
rect 5441 35 5507 38
rect 23933 35 23999 38
rect 36997 98 37063 101
rect 54017 98 54083 101
rect 36997 96 54083 98
rect 36997 40 37002 96
rect 37058 40 54022 96
rect 54078 40 54083 96
rect 36997 38 54083 40
rect 36997 35 37063 38
rect 54017 35 54083 38
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 -7066 -8106 711002
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 -6106 -7146 710042
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 -5146 -6186 709082
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 -4186 -5226 708122
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 -3226 -4266 707162
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 -2266 -3306 706202
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 694354 -2346 705242
rect 582294 705798 582914 711590
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 582294 705562 582326 705798
rect 582562 705562 582646 705798
rect 582882 705562 582914 705798
rect 582294 705478 582914 705562
rect 582294 705242 582326 705478
rect 582562 705242 582646 705478
rect 582882 705242 582914 705478
rect -2966 694118 -2934 694354
rect -2698 694118 -2614 694354
rect -2378 694118 -2346 694354
rect -2966 694034 -2346 694118
rect -2966 693798 -2934 694034
rect -2698 693798 -2614 694034
rect -2378 693798 -2346 694034
rect -2966 658354 -2346 693798
rect -2966 658118 -2934 658354
rect -2698 658118 -2614 658354
rect -2378 658118 -2346 658354
rect -2966 658034 -2346 658118
rect -2966 657798 -2934 658034
rect -2698 657798 -2614 658034
rect -2378 657798 -2346 658034
rect -2966 622354 -2346 657798
rect -2966 622118 -2934 622354
rect -2698 622118 -2614 622354
rect -2378 622118 -2346 622354
rect -2966 622034 -2346 622118
rect -2966 621798 -2934 622034
rect -2698 621798 -2614 622034
rect -2378 621798 -2346 622034
rect -2966 586354 -2346 621798
rect -2966 586118 -2934 586354
rect -2698 586118 -2614 586354
rect -2378 586118 -2346 586354
rect -2966 586034 -2346 586118
rect -2966 585798 -2934 586034
rect -2698 585798 -2614 586034
rect -2378 585798 -2346 586034
rect -2966 550354 -2346 585798
rect -2966 550118 -2934 550354
rect -2698 550118 -2614 550354
rect -2378 550118 -2346 550354
rect -2966 550034 -2346 550118
rect -2966 549798 -2934 550034
rect -2698 549798 -2614 550034
rect -2378 549798 -2346 550034
rect -2966 514354 -2346 549798
rect -2966 514118 -2934 514354
rect -2698 514118 -2614 514354
rect -2378 514118 -2346 514354
rect -2966 514034 -2346 514118
rect -2966 513798 -2934 514034
rect -2698 513798 -2614 514034
rect -2378 513798 -2346 514034
rect -2966 478354 -2346 513798
rect -2966 478118 -2934 478354
rect -2698 478118 -2614 478354
rect -2378 478118 -2346 478354
rect -2966 478034 -2346 478118
rect -2966 477798 -2934 478034
rect -2698 477798 -2614 478034
rect -2378 477798 -2346 478034
rect -2966 442354 -2346 477798
rect -2966 442118 -2934 442354
rect -2698 442118 -2614 442354
rect -2378 442118 -2346 442354
rect -2966 442034 -2346 442118
rect -2966 441798 -2934 442034
rect -2698 441798 -2614 442034
rect -2378 441798 -2346 442034
rect -2966 406354 -2346 441798
rect -2966 406118 -2934 406354
rect -2698 406118 -2614 406354
rect -2378 406118 -2346 406354
rect -2966 406034 -2346 406118
rect -2966 405798 -2934 406034
rect -2698 405798 -2614 406034
rect -2378 405798 -2346 406034
rect -2966 370354 -2346 405798
rect -2966 370118 -2934 370354
rect -2698 370118 -2614 370354
rect -2378 370118 -2346 370354
rect -2966 370034 -2346 370118
rect -2966 369798 -2934 370034
rect -2698 369798 -2614 370034
rect -2378 369798 -2346 370034
rect -2966 334354 -2346 369798
rect -2966 334118 -2934 334354
rect -2698 334118 -2614 334354
rect -2378 334118 -2346 334354
rect -2966 334034 -2346 334118
rect -2966 333798 -2934 334034
rect -2698 333798 -2614 334034
rect -2378 333798 -2346 334034
rect -2966 298354 -2346 333798
rect -2966 298118 -2934 298354
rect -2698 298118 -2614 298354
rect -2378 298118 -2346 298354
rect -2966 298034 -2346 298118
rect -2966 297798 -2934 298034
rect -2698 297798 -2614 298034
rect -2378 297798 -2346 298034
rect -2966 262354 -2346 297798
rect -2966 262118 -2934 262354
rect -2698 262118 -2614 262354
rect -2378 262118 -2346 262354
rect -2966 262034 -2346 262118
rect -2966 261798 -2934 262034
rect -2698 261798 -2614 262034
rect -2378 261798 -2346 262034
rect -2966 226354 -2346 261798
rect -2966 226118 -2934 226354
rect -2698 226118 -2614 226354
rect -2378 226118 -2346 226354
rect -2966 226034 -2346 226118
rect -2966 225798 -2934 226034
rect -2698 225798 -2614 226034
rect -2378 225798 -2346 226034
rect -2966 190354 -2346 225798
rect -2966 190118 -2934 190354
rect -2698 190118 -2614 190354
rect -2378 190118 -2346 190354
rect -2966 190034 -2346 190118
rect -2966 189798 -2934 190034
rect -2698 189798 -2614 190034
rect -2378 189798 -2346 190034
rect -2966 154354 -2346 189798
rect -2966 154118 -2934 154354
rect -2698 154118 -2614 154354
rect -2378 154118 -2346 154354
rect -2966 154034 -2346 154118
rect -2966 153798 -2934 154034
rect -2698 153798 -2614 154034
rect -2378 153798 -2346 154034
rect -2966 118354 -2346 153798
rect -2966 118118 -2934 118354
rect -2698 118118 -2614 118354
rect -2378 118118 -2346 118354
rect -2966 118034 -2346 118118
rect -2966 117798 -2934 118034
rect -2698 117798 -2614 118034
rect -2378 117798 -2346 118034
rect -2966 82354 -2346 117798
rect -2966 82118 -2934 82354
rect -2698 82118 -2614 82354
rect -2378 82118 -2346 82354
rect -2966 82034 -2346 82118
rect -2966 81798 -2934 82034
rect -2698 81798 -2614 82034
rect -2378 81798 -2346 82034
rect -2966 46354 -2346 81798
rect -2966 46118 -2934 46354
rect -2698 46118 -2614 46354
rect -2378 46118 -2346 46354
rect -2966 46034 -2346 46118
rect -2966 45798 -2934 46034
rect -2698 45798 -2614 46034
rect -2378 45798 -2346 46034
rect -2966 10354 -2346 45798
rect -2966 10118 -2934 10354
rect -2698 10118 -2614 10354
rect -2378 10118 -2346 10354
rect -2966 10034 -2346 10118
rect -2966 9798 -2934 10034
rect -2698 9798 -2614 10034
rect -2378 9798 -2346 10034
rect -2966 -1306 -2346 9798
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 689854 -1386 704282
rect 582294 694354 582914 705242
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 23794 694118 23826 694354
rect 24062 694118 24146 694354
rect 24382 694118 24414 694354
rect 23794 694034 24414 694118
rect 23794 693798 23826 694034
rect 24062 693798 24146 694034
rect 24382 693798 24414 694034
rect 59794 694118 59826 694354
rect 60062 694118 60146 694354
rect 60382 694118 60414 694354
rect 59794 694034 60414 694118
rect 59794 693798 59826 694034
rect 60062 693798 60146 694034
rect 60382 693798 60414 694034
rect 95794 694118 95826 694354
rect 96062 694118 96146 694354
rect 96382 694118 96414 694354
rect 95794 694034 96414 694118
rect 95794 693798 95826 694034
rect 96062 693798 96146 694034
rect 96382 693798 96414 694034
rect 131794 694118 131826 694354
rect 132062 694118 132146 694354
rect 132382 694118 132414 694354
rect 131794 694034 132414 694118
rect 131794 693798 131826 694034
rect 132062 693798 132146 694034
rect 132382 693798 132414 694034
rect 167794 694118 167826 694354
rect 168062 694118 168146 694354
rect 168382 694118 168414 694354
rect 167794 694034 168414 694118
rect 167794 693798 167826 694034
rect 168062 693798 168146 694034
rect 168382 693798 168414 694034
rect 203794 694118 203826 694354
rect 204062 694118 204146 694354
rect 204382 694118 204414 694354
rect 203794 694034 204414 694118
rect 203794 693798 203826 694034
rect 204062 693798 204146 694034
rect 204382 693798 204414 694034
rect 239794 694118 239826 694354
rect 240062 694118 240146 694354
rect 240382 694118 240414 694354
rect 239794 694034 240414 694118
rect 239794 693798 239826 694034
rect 240062 693798 240146 694034
rect 240382 693798 240414 694034
rect 275794 694118 275826 694354
rect 276062 694118 276146 694354
rect 276382 694118 276414 694354
rect 275794 694034 276414 694118
rect 275794 693798 275826 694034
rect 276062 693798 276146 694034
rect 276382 693798 276414 694034
rect 311794 694118 311826 694354
rect 312062 694118 312146 694354
rect 312382 694118 312414 694354
rect 311794 694034 312414 694118
rect 311794 693798 311826 694034
rect 312062 693798 312146 694034
rect 312382 693798 312414 694034
rect 347794 694118 347826 694354
rect 348062 694118 348146 694354
rect 348382 694118 348414 694354
rect 347794 694034 348414 694118
rect 347794 693798 347826 694034
rect 348062 693798 348146 694034
rect 348382 693798 348414 694034
rect 383794 694118 383826 694354
rect 384062 694118 384146 694354
rect 384382 694118 384414 694354
rect 383794 694034 384414 694118
rect 383794 693798 383826 694034
rect 384062 693798 384146 694034
rect 384382 693798 384414 694034
rect 419794 694118 419826 694354
rect 420062 694118 420146 694354
rect 420382 694118 420414 694354
rect 419794 694034 420414 694118
rect 419794 693798 419826 694034
rect 420062 693798 420146 694034
rect 420382 693798 420414 694034
rect 455794 694118 455826 694354
rect 456062 694118 456146 694354
rect 456382 694118 456414 694354
rect 455794 694034 456414 694118
rect 455794 693798 455826 694034
rect 456062 693798 456146 694034
rect 456382 693798 456414 694034
rect 491794 694118 491826 694354
rect 492062 694118 492146 694354
rect 492382 694118 492414 694354
rect 491794 694034 492414 694118
rect 491794 693798 491826 694034
rect 492062 693798 492146 694034
rect 492382 693798 492414 694034
rect 527794 694118 527826 694354
rect 528062 694118 528146 694354
rect 528382 694118 528414 694354
rect 527794 694034 528414 694118
rect 527794 693798 527826 694034
rect 528062 693798 528146 694034
rect 528382 693798 528414 694034
rect 563794 694118 563826 694354
rect 564062 694118 564146 694354
rect 564382 694118 564414 694354
rect 563794 694034 564414 694118
rect 563794 693798 563826 694034
rect 564062 693798 564146 694034
rect 564382 693798 564414 694034
rect 582294 694118 582326 694354
rect 582562 694118 582646 694354
rect 582882 694118 582914 694354
rect 582294 694034 582914 694118
rect 582294 693798 582326 694034
rect 582562 693798 582646 694034
rect 582882 693798 582914 694034
rect -2006 689618 -1974 689854
rect -1738 689618 -1654 689854
rect -1418 689618 -1386 689854
rect -2006 689534 -1386 689618
rect -2006 689298 -1974 689534
rect -1738 689298 -1654 689534
rect -1418 689298 -1386 689534
rect 5794 689618 5826 689854
rect 6062 689618 6146 689854
rect 6382 689618 6414 689854
rect 5794 689534 6414 689618
rect 5794 689298 5826 689534
rect 6062 689298 6146 689534
rect 6382 689298 6414 689534
rect 41794 689618 41826 689854
rect 42062 689618 42146 689854
rect 42382 689618 42414 689854
rect 41794 689534 42414 689618
rect 41794 689298 41826 689534
rect 42062 689298 42146 689534
rect 42382 689298 42414 689534
rect 77794 689618 77826 689854
rect 78062 689618 78146 689854
rect 78382 689618 78414 689854
rect 77794 689534 78414 689618
rect 77794 689298 77826 689534
rect 78062 689298 78146 689534
rect 78382 689298 78414 689534
rect 113794 689618 113826 689854
rect 114062 689618 114146 689854
rect 114382 689618 114414 689854
rect 113794 689534 114414 689618
rect 113794 689298 113826 689534
rect 114062 689298 114146 689534
rect 114382 689298 114414 689534
rect 149794 689618 149826 689854
rect 150062 689618 150146 689854
rect 150382 689618 150414 689854
rect 149794 689534 150414 689618
rect 149794 689298 149826 689534
rect 150062 689298 150146 689534
rect 150382 689298 150414 689534
rect 185794 689618 185826 689854
rect 186062 689618 186146 689854
rect 186382 689618 186414 689854
rect 185794 689534 186414 689618
rect 185794 689298 185826 689534
rect 186062 689298 186146 689534
rect 186382 689298 186414 689534
rect 221794 689618 221826 689854
rect 222062 689618 222146 689854
rect 222382 689618 222414 689854
rect 221794 689534 222414 689618
rect 221794 689298 221826 689534
rect 222062 689298 222146 689534
rect 222382 689298 222414 689534
rect 257794 689618 257826 689854
rect 258062 689618 258146 689854
rect 258382 689618 258414 689854
rect 257794 689534 258414 689618
rect 257794 689298 257826 689534
rect 258062 689298 258146 689534
rect 258382 689298 258414 689534
rect 293794 689618 293826 689854
rect 294062 689618 294146 689854
rect 294382 689618 294414 689854
rect 293794 689534 294414 689618
rect 293794 689298 293826 689534
rect 294062 689298 294146 689534
rect 294382 689298 294414 689534
rect 329794 689618 329826 689854
rect 330062 689618 330146 689854
rect 330382 689618 330414 689854
rect 329794 689534 330414 689618
rect 329794 689298 329826 689534
rect 330062 689298 330146 689534
rect 330382 689298 330414 689534
rect 365794 689618 365826 689854
rect 366062 689618 366146 689854
rect 366382 689618 366414 689854
rect 365794 689534 366414 689618
rect 365794 689298 365826 689534
rect 366062 689298 366146 689534
rect 366382 689298 366414 689534
rect 401794 689618 401826 689854
rect 402062 689618 402146 689854
rect 402382 689618 402414 689854
rect 401794 689534 402414 689618
rect 401794 689298 401826 689534
rect 402062 689298 402146 689534
rect 402382 689298 402414 689534
rect 437794 689618 437826 689854
rect 438062 689618 438146 689854
rect 438382 689618 438414 689854
rect 437794 689534 438414 689618
rect 437794 689298 437826 689534
rect 438062 689298 438146 689534
rect 438382 689298 438414 689534
rect 473794 689618 473826 689854
rect 474062 689618 474146 689854
rect 474382 689618 474414 689854
rect 473794 689534 474414 689618
rect 473794 689298 473826 689534
rect 474062 689298 474146 689534
rect 474382 689298 474414 689534
rect 509794 689618 509826 689854
rect 510062 689618 510146 689854
rect 510382 689618 510414 689854
rect 509794 689534 510414 689618
rect 509794 689298 509826 689534
rect 510062 689298 510146 689534
rect 510382 689298 510414 689534
rect 545794 689618 545826 689854
rect 546062 689618 546146 689854
rect 546382 689618 546414 689854
rect 545794 689534 546414 689618
rect 545794 689298 545826 689534
rect 546062 689298 546146 689534
rect 546382 689298 546414 689534
rect -2006 653854 -1386 689298
rect 582294 658354 582914 693798
rect 13166 658118 13198 658354
rect 13434 658118 13518 658354
rect 13754 658118 13786 658354
rect 13166 658034 13786 658118
rect 13166 657798 13198 658034
rect 13434 657798 13518 658034
rect 13754 657798 13786 658034
rect 167794 658118 167826 658354
rect 168062 658118 168146 658354
rect 168382 658118 168414 658354
rect 167794 658034 168414 658118
rect 167794 657798 167826 658034
rect 168062 657798 168146 658034
rect 168382 657798 168414 658034
rect 291558 658118 291590 658354
rect 291826 658118 291910 658354
rect 292146 658118 292178 658354
rect 291558 658034 292178 658118
rect 291558 657798 291590 658034
rect 291826 657798 291910 658034
rect 292146 657798 292178 658034
rect 419794 658118 419826 658354
rect 420062 658118 420146 658354
rect 420382 658118 420414 658354
rect 419794 658034 420414 658118
rect 419794 657798 419826 658034
rect 420062 657798 420146 658034
rect 420382 657798 420414 658034
rect 563794 658118 563826 658354
rect 564062 658118 564146 658354
rect 564382 658118 564414 658354
rect 563794 658034 564414 658118
rect 563794 657798 563826 658034
rect 564062 657798 564146 658034
rect 564382 657798 564414 658034
rect 582294 658118 582326 658354
rect 582562 658118 582646 658354
rect 582882 658118 582914 658354
rect 582294 658034 582914 658118
rect 582294 657798 582326 658034
rect 582562 657798 582646 658034
rect 582882 657798 582914 658034
rect -2006 653618 -1974 653854
rect -1738 653618 -1654 653854
rect -1418 653618 -1386 653854
rect -2006 653534 -1386 653618
rect -2006 653298 -1974 653534
rect -1738 653298 -1654 653534
rect -1418 653298 -1386 653534
rect 5794 653618 5826 653854
rect 6062 653618 6146 653854
rect 6382 653618 6414 653854
rect 5794 653534 6414 653618
rect 5794 653298 5826 653534
rect 6062 653298 6146 653534
rect 6382 653298 6414 653534
rect 173062 653618 173094 653854
rect 173330 653618 173414 653854
rect 173650 653618 173682 653854
rect 173062 653534 173682 653618
rect 173062 653298 173094 653534
rect 173330 653298 173414 653534
rect 173650 653298 173682 653534
rect 293794 653618 293826 653854
rect 294062 653618 294146 653854
rect 294382 653618 294414 653854
rect 293794 653534 294414 653618
rect 293794 653298 293826 653534
rect 294062 653298 294146 653534
rect 294382 653298 294414 653534
rect 401794 653618 401826 653854
rect 402062 653618 402146 653854
rect 402382 653618 402414 653854
rect 401794 653534 402414 653618
rect 401794 653298 401826 653534
rect 402062 653298 402146 653534
rect 402382 653298 402414 653534
rect 570318 653618 570350 653854
rect 570586 653618 570670 653854
rect 570906 653618 570938 653854
rect 570318 653534 570938 653618
rect 570318 653298 570350 653534
rect 570586 653298 570670 653534
rect 570906 653298 570938 653534
rect -2006 617854 -1386 653298
rect 582294 622354 582914 657798
rect 13166 622118 13198 622354
rect 13434 622118 13518 622354
rect 13754 622118 13786 622354
rect 13166 622034 13786 622118
rect 13166 621798 13198 622034
rect 13434 621798 13518 622034
rect 13754 621798 13786 622034
rect 167794 622118 167826 622354
rect 168062 622118 168146 622354
rect 168382 622118 168414 622354
rect 167794 622034 168414 622118
rect 167794 621798 167826 622034
rect 168062 621798 168146 622034
rect 168382 621798 168414 622034
rect 291558 622118 291590 622354
rect 291826 622118 291910 622354
rect 292146 622118 292178 622354
rect 291558 622034 292178 622118
rect 291558 621798 291590 622034
rect 291826 621798 291910 622034
rect 292146 621798 292178 622034
rect 419794 622118 419826 622354
rect 420062 622118 420146 622354
rect 420382 622118 420414 622354
rect 419794 622034 420414 622118
rect 419794 621798 419826 622034
rect 420062 621798 420146 622034
rect 420382 621798 420414 622034
rect 563794 622118 563826 622354
rect 564062 622118 564146 622354
rect 564382 622118 564414 622354
rect 563794 622034 564414 622118
rect 563794 621798 563826 622034
rect 564062 621798 564146 622034
rect 564382 621798 564414 622034
rect 582294 622118 582326 622354
rect 582562 622118 582646 622354
rect 582882 622118 582914 622354
rect 582294 622034 582914 622118
rect 582294 621798 582326 622034
rect 582562 621798 582646 622034
rect 582882 621798 582914 622034
rect -2006 617618 -1974 617854
rect -1738 617618 -1654 617854
rect -1418 617618 -1386 617854
rect -2006 617534 -1386 617618
rect -2006 617298 -1974 617534
rect -1738 617298 -1654 617534
rect -1418 617298 -1386 617534
rect 5794 617618 5826 617854
rect 6062 617618 6146 617854
rect 6382 617618 6414 617854
rect 5794 617534 6414 617618
rect 5794 617298 5826 617534
rect 6062 617298 6146 617534
rect 6382 617298 6414 617534
rect 173062 617618 173094 617854
rect 173330 617618 173414 617854
rect 173650 617618 173682 617854
rect 173062 617534 173682 617618
rect 173062 617298 173094 617534
rect 173330 617298 173414 617534
rect 173650 617298 173682 617534
rect 293794 617618 293826 617854
rect 294062 617618 294146 617854
rect 294382 617618 294414 617854
rect 293794 617534 294414 617618
rect 293794 617298 293826 617534
rect 294062 617298 294146 617534
rect 294382 617298 294414 617534
rect 401794 617618 401826 617854
rect 402062 617618 402146 617854
rect 402382 617618 402414 617854
rect 401794 617534 402414 617618
rect 401794 617298 401826 617534
rect 402062 617298 402146 617534
rect 402382 617298 402414 617534
rect 570318 617618 570350 617854
rect 570586 617618 570670 617854
rect 570906 617618 570938 617854
rect 570318 617534 570938 617618
rect 570318 617298 570350 617534
rect 570586 617298 570670 617534
rect 570906 617298 570938 617534
rect -2006 581854 -1386 617298
rect 582294 586354 582914 621798
rect 23794 586118 23826 586354
rect 24062 586118 24146 586354
rect 24382 586118 24414 586354
rect 23794 586034 24414 586118
rect 23794 585798 23826 586034
rect 24062 585798 24146 586034
rect 24382 585798 24414 586034
rect 59794 586118 59826 586354
rect 60062 586118 60146 586354
rect 60382 586118 60414 586354
rect 59794 586034 60414 586118
rect 59794 585798 59826 586034
rect 60062 585798 60146 586034
rect 60382 585798 60414 586034
rect 95794 586118 95826 586354
rect 96062 586118 96146 586354
rect 96382 586118 96414 586354
rect 95794 586034 96414 586118
rect 95794 585798 95826 586034
rect 96062 585798 96146 586034
rect 96382 585798 96414 586034
rect 131794 586118 131826 586354
rect 132062 586118 132146 586354
rect 132382 586118 132414 586354
rect 131794 586034 132414 586118
rect 131794 585798 131826 586034
rect 132062 585798 132146 586034
rect 132382 585798 132414 586034
rect 167794 586118 167826 586354
rect 168062 586118 168146 586354
rect 168382 586118 168414 586354
rect 167794 586034 168414 586118
rect 167794 585798 167826 586034
rect 168062 585798 168146 586034
rect 168382 585798 168414 586034
rect 203794 586118 203826 586354
rect 204062 586118 204146 586354
rect 204382 586118 204414 586354
rect 203794 586034 204414 586118
rect 203794 585798 203826 586034
rect 204062 585798 204146 586034
rect 204382 585798 204414 586034
rect 239794 586118 239826 586354
rect 240062 586118 240146 586354
rect 240382 586118 240414 586354
rect 239794 586034 240414 586118
rect 239794 585798 239826 586034
rect 240062 585798 240146 586034
rect 240382 585798 240414 586034
rect 275794 586118 275826 586354
rect 276062 586118 276146 586354
rect 276382 586118 276414 586354
rect 275794 586034 276414 586118
rect 275794 585798 275826 586034
rect 276062 585798 276146 586034
rect 276382 585798 276414 586034
rect 311794 586118 311826 586354
rect 312062 586118 312146 586354
rect 312382 586118 312414 586354
rect 311794 586034 312414 586118
rect 311794 585798 311826 586034
rect 312062 585798 312146 586034
rect 312382 585798 312414 586034
rect 347794 586118 347826 586354
rect 348062 586118 348146 586354
rect 348382 586118 348414 586354
rect 347794 586034 348414 586118
rect 347794 585798 347826 586034
rect 348062 585798 348146 586034
rect 348382 585798 348414 586034
rect 383794 586118 383826 586354
rect 384062 586118 384146 586354
rect 384382 586118 384414 586354
rect 383794 586034 384414 586118
rect 383794 585798 383826 586034
rect 384062 585798 384146 586034
rect 384382 585798 384414 586034
rect 419794 586118 419826 586354
rect 420062 586118 420146 586354
rect 420382 586118 420414 586354
rect 419794 586034 420414 586118
rect 419794 585798 419826 586034
rect 420062 585798 420146 586034
rect 420382 585798 420414 586034
rect 455794 586118 455826 586354
rect 456062 586118 456146 586354
rect 456382 586118 456414 586354
rect 455794 586034 456414 586118
rect 455794 585798 455826 586034
rect 456062 585798 456146 586034
rect 456382 585798 456414 586034
rect 491794 586118 491826 586354
rect 492062 586118 492146 586354
rect 492382 586118 492414 586354
rect 491794 586034 492414 586118
rect 491794 585798 491826 586034
rect 492062 585798 492146 586034
rect 492382 585798 492414 586034
rect 527794 586118 527826 586354
rect 528062 586118 528146 586354
rect 528382 586118 528414 586354
rect 527794 586034 528414 586118
rect 527794 585798 527826 586034
rect 528062 585798 528146 586034
rect 528382 585798 528414 586034
rect 563794 586118 563826 586354
rect 564062 586118 564146 586354
rect 564382 586118 564414 586354
rect 563794 586034 564414 586118
rect 563794 585798 563826 586034
rect 564062 585798 564146 586034
rect 564382 585798 564414 586034
rect 582294 586118 582326 586354
rect 582562 586118 582646 586354
rect 582882 586118 582914 586354
rect 582294 586034 582914 586118
rect 582294 585798 582326 586034
rect 582562 585798 582646 586034
rect 582882 585798 582914 586034
rect -2006 581618 -1974 581854
rect -1738 581618 -1654 581854
rect -1418 581618 -1386 581854
rect -2006 581534 -1386 581618
rect -2006 581298 -1974 581534
rect -1738 581298 -1654 581534
rect -1418 581298 -1386 581534
rect 5794 581618 5826 581854
rect 6062 581618 6146 581854
rect 6382 581618 6414 581854
rect 5794 581534 6414 581618
rect 5794 581298 5826 581534
rect 6062 581298 6146 581534
rect 6382 581298 6414 581534
rect 41794 581618 41826 581854
rect 42062 581618 42146 581854
rect 42382 581618 42414 581854
rect 41794 581534 42414 581618
rect 41794 581298 41826 581534
rect 42062 581298 42146 581534
rect 42382 581298 42414 581534
rect 77794 581618 77826 581854
rect 78062 581618 78146 581854
rect 78382 581618 78414 581854
rect 77794 581534 78414 581618
rect 77794 581298 77826 581534
rect 78062 581298 78146 581534
rect 78382 581298 78414 581534
rect 113794 581618 113826 581854
rect 114062 581618 114146 581854
rect 114382 581618 114414 581854
rect 113794 581534 114414 581618
rect 113794 581298 113826 581534
rect 114062 581298 114146 581534
rect 114382 581298 114414 581534
rect 149794 581618 149826 581854
rect 150062 581618 150146 581854
rect 150382 581618 150414 581854
rect 149794 581534 150414 581618
rect 149794 581298 149826 581534
rect 150062 581298 150146 581534
rect 150382 581298 150414 581534
rect 185794 581618 185826 581854
rect 186062 581618 186146 581854
rect 186382 581618 186414 581854
rect 185794 581534 186414 581618
rect 185794 581298 185826 581534
rect 186062 581298 186146 581534
rect 186382 581298 186414 581534
rect 221794 581618 221826 581854
rect 222062 581618 222146 581854
rect 222382 581618 222414 581854
rect 221794 581534 222414 581618
rect 221794 581298 221826 581534
rect 222062 581298 222146 581534
rect 222382 581298 222414 581534
rect 257794 581618 257826 581854
rect 258062 581618 258146 581854
rect 258382 581618 258414 581854
rect 257794 581534 258414 581618
rect 257794 581298 257826 581534
rect 258062 581298 258146 581534
rect 258382 581298 258414 581534
rect 293794 581618 293826 581854
rect 294062 581618 294146 581854
rect 294382 581618 294414 581854
rect 293794 581534 294414 581618
rect 293794 581298 293826 581534
rect 294062 581298 294146 581534
rect 294382 581298 294414 581534
rect 329794 581618 329826 581854
rect 330062 581618 330146 581854
rect 330382 581618 330414 581854
rect 329794 581534 330414 581618
rect 329794 581298 329826 581534
rect 330062 581298 330146 581534
rect 330382 581298 330414 581534
rect 365794 581618 365826 581854
rect 366062 581618 366146 581854
rect 366382 581618 366414 581854
rect 365794 581534 366414 581618
rect 365794 581298 365826 581534
rect 366062 581298 366146 581534
rect 366382 581298 366414 581534
rect 401794 581618 401826 581854
rect 402062 581618 402146 581854
rect 402382 581618 402414 581854
rect 401794 581534 402414 581618
rect 401794 581298 401826 581534
rect 402062 581298 402146 581534
rect 402382 581298 402414 581534
rect 437794 581618 437826 581854
rect 438062 581618 438146 581854
rect 438382 581618 438414 581854
rect 437794 581534 438414 581618
rect 437794 581298 437826 581534
rect 438062 581298 438146 581534
rect 438382 581298 438414 581534
rect 473794 581618 473826 581854
rect 474062 581618 474146 581854
rect 474382 581618 474414 581854
rect 473794 581534 474414 581618
rect 473794 581298 473826 581534
rect 474062 581298 474146 581534
rect 474382 581298 474414 581534
rect 509794 581618 509826 581854
rect 510062 581618 510146 581854
rect 510382 581618 510414 581854
rect 509794 581534 510414 581618
rect 509794 581298 509826 581534
rect 510062 581298 510146 581534
rect 510382 581298 510414 581534
rect 545794 581618 545826 581854
rect 546062 581618 546146 581854
rect 546382 581618 546414 581854
rect 545794 581534 546414 581618
rect 545794 581298 545826 581534
rect 546062 581298 546146 581534
rect 546382 581298 546414 581534
rect -2006 545854 -1386 581298
rect 582294 550354 582914 585798
rect 13166 550118 13198 550354
rect 13434 550118 13518 550354
rect 13754 550118 13786 550354
rect 13166 550034 13786 550118
rect 13166 549798 13198 550034
rect 13434 549798 13518 550034
rect 13754 549798 13786 550034
rect 167794 550118 167826 550354
rect 168062 550118 168146 550354
rect 168382 550118 168414 550354
rect 167794 550034 168414 550118
rect 167794 549798 167826 550034
rect 168062 549798 168146 550034
rect 168382 549798 168414 550034
rect 203794 550118 203826 550354
rect 204062 550118 204146 550354
rect 204382 550118 204414 550354
rect 203794 550034 204414 550118
rect 203794 549798 203826 550034
rect 204062 549798 204146 550034
rect 204382 549798 204414 550034
rect 239794 550118 239826 550354
rect 240062 550118 240146 550354
rect 240382 550118 240414 550354
rect 239794 550034 240414 550118
rect 239794 549798 239826 550034
rect 240062 549798 240146 550034
rect 240382 549798 240414 550034
rect 275794 550118 275826 550354
rect 276062 550118 276146 550354
rect 276382 550118 276414 550354
rect 275794 550034 276414 550118
rect 275794 549798 275826 550034
rect 276062 549798 276146 550034
rect 276382 549798 276414 550034
rect 311794 550118 311826 550354
rect 312062 550118 312146 550354
rect 312382 550118 312414 550354
rect 311794 550034 312414 550118
rect 311794 549798 311826 550034
rect 312062 549798 312146 550034
rect 312382 549798 312414 550034
rect 347794 550118 347826 550354
rect 348062 550118 348146 550354
rect 348382 550118 348414 550354
rect 347794 550034 348414 550118
rect 347794 549798 347826 550034
rect 348062 549798 348146 550034
rect 348382 549798 348414 550034
rect 383794 550118 383826 550354
rect 384062 550118 384146 550354
rect 384382 550118 384414 550354
rect 383794 550034 384414 550118
rect 383794 549798 383826 550034
rect 384062 549798 384146 550034
rect 384382 549798 384414 550034
rect 419794 550118 419826 550354
rect 420062 550118 420146 550354
rect 420382 550118 420414 550354
rect 419794 550034 420414 550118
rect 419794 549798 419826 550034
rect 420062 549798 420146 550034
rect 420382 549798 420414 550034
rect 563794 550118 563826 550354
rect 564062 550118 564146 550354
rect 564382 550118 564414 550354
rect 563794 550034 564414 550118
rect 563794 549798 563826 550034
rect 564062 549798 564146 550034
rect 564382 549798 564414 550034
rect 582294 550118 582326 550354
rect 582562 550118 582646 550354
rect 582882 550118 582914 550354
rect 582294 550034 582914 550118
rect 582294 549798 582326 550034
rect 582562 549798 582646 550034
rect 582882 549798 582914 550034
rect -2006 545618 -1974 545854
rect -1738 545618 -1654 545854
rect -1418 545618 -1386 545854
rect -2006 545534 -1386 545618
rect -2006 545298 -1974 545534
rect -1738 545298 -1654 545534
rect -1418 545298 -1386 545534
rect 5794 545618 5826 545854
rect 6062 545618 6146 545854
rect 6382 545618 6414 545854
rect 5794 545534 6414 545618
rect 5794 545298 5826 545534
rect 6062 545298 6146 545534
rect 6382 545298 6414 545534
rect 185794 545618 185826 545854
rect 186062 545618 186146 545854
rect 186382 545618 186414 545854
rect 185794 545534 186414 545618
rect 185794 545298 185826 545534
rect 186062 545298 186146 545534
rect 186382 545298 186414 545534
rect 221794 545618 221826 545854
rect 222062 545618 222146 545854
rect 222382 545618 222414 545854
rect 221794 545534 222414 545618
rect 221794 545298 221826 545534
rect 222062 545298 222146 545534
rect 222382 545298 222414 545534
rect 257794 545618 257826 545854
rect 258062 545618 258146 545854
rect 258382 545618 258414 545854
rect 257794 545534 258414 545618
rect 257794 545298 257826 545534
rect 258062 545298 258146 545534
rect 258382 545298 258414 545534
rect 293794 545618 293826 545854
rect 294062 545618 294146 545854
rect 294382 545618 294414 545854
rect 293794 545534 294414 545618
rect 293794 545298 293826 545534
rect 294062 545298 294146 545534
rect 294382 545298 294414 545534
rect 329794 545618 329826 545854
rect 330062 545618 330146 545854
rect 330382 545618 330414 545854
rect 329794 545534 330414 545618
rect 329794 545298 329826 545534
rect 330062 545298 330146 545534
rect 330382 545298 330414 545534
rect 365794 545618 365826 545854
rect 366062 545618 366146 545854
rect 366382 545618 366414 545854
rect 365794 545534 366414 545618
rect 365794 545298 365826 545534
rect 366062 545298 366146 545534
rect 366382 545298 366414 545534
rect 401794 545618 401826 545854
rect 402062 545618 402146 545854
rect 402382 545618 402414 545854
rect 401794 545534 402414 545618
rect 401794 545298 401826 545534
rect 402062 545298 402146 545534
rect 402382 545298 402414 545534
rect 570318 545618 570350 545854
rect 570586 545618 570670 545854
rect 570906 545618 570938 545854
rect 570318 545534 570938 545618
rect 570318 545298 570350 545534
rect 570586 545298 570670 545534
rect 570906 545298 570938 545534
rect -2006 509854 -1386 545298
rect 582294 514354 582914 549798
rect 13166 514118 13198 514354
rect 13434 514118 13518 514354
rect 13754 514118 13786 514354
rect 13166 514034 13786 514118
rect 13166 513798 13198 514034
rect 13434 513798 13518 514034
rect 13754 513798 13786 514034
rect 167794 514118 167826 514354
rect 168062 514118 168146 514354
rect 168382 514118 168414 514354
rect 167794 514034 168414 514118
rect 167794 513798 167826 514034
rect 168062 513798 168146 514034
rect 168382 513798 168414 514034
rect 203794 514118 203826 514354
rect 204062 514118 204146 514354
rect 204382 514118 204414 514354
rect 203794 514034 204414 514118
rect 203794 513798 203826 514034
rect 204062 513798 204146 514034
rect 204382 513798 204414 514034
rect 239794 514118 239826 514354
rect 240062 514118 240146 514354
rect 240382 514118 240414 514354
rect 239794 514034 240414 514118
rect 239794 513798 239826 514034
rect 240062 513798 240146 514034
rect 240382 513798 240414 514034
rect 275794 514118 275826 514354
rect 276062 514118 276146 514354
rect 276382 514118 276414 514354
rect 275794 514034 276414 514118
rect 275794 513798 275826 514034
rect 276062 513798 276146 514034
rect 276382 513798 276414 514034
rect 311794 514118 311826 514354
rect 312062 514118 312146 514354
rect 312382 514118 312414 514354
rect 311794 514034 312414 514118
rect 311794 513798 311826 514034
rect 312062 513798 312146 514034
rect 312382 513798 312414 514034
rect 347794 514118 347826 514354
rect 348062 514118 348146 514354
rect 348382 514118 348414 514354
rect 347794 514034 348414 514118
rect 347794 513798 347826 514034
rect 348062 513798 348146 514034
rect 348382 513798 348414 514034
rect 383794 514118 383826 514354
rect 384062 514118 384146 514354
rect 384382 514118 384414 514354
rect 383794 514034 384414 514118
rect 383794 513798 383826 514034
rect 384062 513798 384146 514034
rect 384382 513798 384414 514034
rect 419794 514118 419826 514354
rect 420062 514118 420146 514354
rect 420382 514118 420414 514354
rect 419794 514034 420414 514118
rect 419794 513798 419826 514034
rect 420062 513798 420146 514034
rect 420382 513798 420414 514034
rect 563794 514118 563826 514354
rect 564062 514118 564146 514354
rect 564382 514118 564414 514354
rect 563794 514034 564414 514118
rect 563794 513798 563826 514034
rect 564062 513798 564146 514034
rect 564382 513798 564414 514034
rect 582294 514118 582326 514354
rect 582562 514118 582646 514354
rect 582882 514118 582914 514354
rect 582294 514034 582914 514118
rect 582294 513798 582326 514034
rect 582562 513798 582646 514034
rect 582882 513798 582914 514034
rect -2006 509618 -1974 509854
rect -1738 509618 -1654 509854
rect -1418 509618 -1386 509854
rect -2006 509534 -1386 509618
rect -2006 509298 -1974 509534
rect -1738 509298 -1654 509534
rect -1418 509298 -1386 509534
rect 5794 509618 5826 509854
rect 6062 509618 6146 509854
rect 6382 509618 6414 509854
rect 5794 509534 6414 509618
rect 5794 509298 5826 509534
rect 6062 509298 6146 509534
rect 6382 509298 6414 509534
rect 185794 509618 185826 509854
rect 186062 509618 186146 509854
rect 186382 509618 186414 509854
rect 185794 509534 186414 509618
rect 185794 509298 185826 509534
rect 186062 509298 186146 509534
rect 186382 509298 186414 509534
rect 221794 509618 221826 509854
rect 222062 509618 222146 509854
rect 222382 509618 222414 509854
rect 221794 509534 222414 509618
rect 221794 509298 221826 509534
rect 222062 509298 222146 509534
rect 222382 509298 222414 509534
rect 257794 509618 257826 509854
rect 258062 509618 258146 509854
rect 258382 509618 258414 509854
rect 257794 509534 258414 509618
rect 257794 509298 257826 509534
rect 258062 509298 258146 509534
rect 258382 509298 258414 509534
rect 293794 509618 293826 509854
rect 294062 509618 294146 509854
rect 294382 509618 294414 509854
rect 293794 509534 294414 509618
rect 293794 509298 293826 509534
rect 294062 509298 294146 509534
rect 294382 509298 294414 509534
rect 329794 509618 329826 509854
rect 330062 509618 330146 509854
rect 330382 509618 330414 509854
rect 329794 509534 330414 509618
rect 329794 509298 329826 509534
rect 330062 509298 330146 509534
rect 330382 509298 330414 509534
rect 365794 509618 365826 509854
rect 366062 509618 366146 509854
rect 366382 509618 366414 509854
rect 365794 509534 366414 509618
rect 365794 509298 365826 509534
rect 366062 509298 366146 509534
rect 366382 509298 366414 509534
rect 401794 509618 401826 509854
rect 402062 509618 402146 509854
rect 402382 509618 402414 509854
rect 401794 509534 402414 509618
rect 401794 509298 401826 509534
rect 402062 509298 402146 509534
rect 402382 509298 402414 509534
rect 570318 509618 570350 509854
rect 570586 509618 570670 509854
rect 570906 509618 570938 509854
rect 570318 509534 570938 509618
rect 570318 509298 570350 509534
rect 570586 509298 570670 509534
rect 570906 509298 570938 509534
rect -2006 473854 -1386 509298
rect 582294 478354 582914 513798
rect 23794 478118 23826 478354
rect 24062 478118 24146 478354
rect 24382 478118 24414 478354
rect 23794 478034 24414 478118
rect 23794 477798 23826 478034
rect 24062 477798 24146 478034
rect 24382 477798 24414 478034
rect 59794 478118 59826 478354
rect 60062 478118 60146 478354
rect 60382 478118 60414 478354
rect 59794 478034 60414 478118
rect 59794 477798 59826 478034
rect 60062 477798 60146 478034
rect 60382 477798 60414 478034
rect 95794 478118 95826 478354
rect 96062 478118 96146 478354
rect 96382 478118 96414 478354
rect 95794 478034 96414 478118
rect 95794 477798 95826 478034
rect 96062 477798 96146 478034
rect 96382 477798 96414 478034
rect 131794 478118 131826 478354
rect 132062 478118 132146 478354
rect 132382 478118 132414 478354
rect 131794 478034 132414 478118
rect 131794 477798 131826 478034
rect 132062 477798 132146 478034
rect 132382 477798 132414 478034
rect 167794 478118 167826 478354
rect 168062 478118 168146 478354
rect 168382 478118 168414 478354
rect 167794 478034 168414 478118
rect 167794 477798 167826 478034
rect 168062 477798 168146 478034
rect 168382 477798 168414 478034
rect 203794 478118 203826 478354
rect 204062 478118 204146 478354
rect 204382 478118 204414 478354
rect 203794 478034 204414 478118
rect 203794 477798 203826 478034
rect 204062 477798 204146 478034
rect 204382 477798 204414 478034
rect 239794 478118 239826 478354
rect 240062 478118 240146 478354
rect 240382 478118 240414 478354
rect 239794 478034 240414 478118
rect 239794 477798 239826 478034
rect 240062 477798 240146 478034
rect 240382 477798 240414 478034
rect 275794 478118 275826 478354
rect 276062 478118 276146 478354
rect 276382 478118 276414 478354
rect 275794 478034 276414 478118
rect 275794 477798 275826 478034
rect 276062 477798 276146 478034
rect 276382 477798 276414 478034
rect 311794 478118 311826 478354
rect 312062 478118 312146 478354
rect 312382 478118 312414 478354
rect 311794 478034 312414 478118
rect 311794 477798 311826 478034
rect 312062 477798 312146 478034
rect 312382 477798 312414 478034
rect 347794 478118 347826 478354
rect 348062 478118 348146 478354
rect 348382 478118 348414 478354
rect 347794 478034 348414 478118
rect 347794 477798 347826 478034
rect 348062 477798 348146 478034
rect 348382 477798 348414 478034
rect 383794 478118 383826 478354
rect 384062 478118 384146 478354
rect 384382 478118 384414 478354
rect 383794 478034 384414 478118
rect 383794 477798 383826 478034
rect 384062 477798 384146 478034
rect 384382 477798 384414 478034
rect 419794 478118 419826 478354
rect 420062 478118 420146 478354
rect 420382 478118 420414 478354
rect 419794 478034 420414 478118
rect 419794 477798 419826 478034
rect 420062 477798 420146 478034
rect 420382 477798 420414 478034
rect 455794 478118 455826 478354
rect 456062 478118 456146 478354
rect 456382 478118 456414 478354
rect 455794 478034 456414 478118
rect 455794 477798 455826 478034
rect 456062 477798 456146 478034
rect 456382 477798 456414 478034
rect 491794 478118 491826 478354
rect 492062 478118 492146 478354
rect 492382 478118 492414 478354
rect 491794 478034 492414 478118
rect 491794 477798 491826 478034
rect 492062 477798 492146 478034
rect 492382 477798 492414 478034
rect 527794 478118 527826 478354
rect 528062 478118 528146 478354
rect 528382 478118 528414 478354
rect 527794 478034 528414 478118
rect 527794 477798 527826 478034
rect 528062 477798 528146 478034
rect 528382 477798 528414 478034
rect 563794 478118 563826 478354
rect 564062 478118 564146 478354
rect 564382 478118 564414 478354
rect 563794 478034 564414 478118
rect 563794 477798 563826 478034
rect 564062 477798 564146 478034
rect 564382 477798 564414 478034
rect 582294 478118 582326 478354
rect 582562 478118 582646 478354
rect 582882 478118 582914 478354
rect 582294 478034 582914 478118
rect 582294 477798 582326 478034
rect 582562 477798 582646 478034
rect 582882 477798 582914 478034
rect -2006 473618 -1974 473854
rect -1738 473618 -1654 473854
rect -1418 473618 -1386 473854
rect -2006 473534 -1386 473618
rect -2006 473298 -1974 473534
rect -1738 473298 -1654 473534
rect -1418 473298 -1386 473534
rect 5794 473618 5826 473854
rect 6062 473618 6146 473854
rect 6382 473618 6414 473854
rect 5794 473534 6414 473618
rect 5794 473298 5826 473534
rect 6062 473298 6146 473534
rect 6382 473298 6414 473534
rect 41794 473618 41826 473854
rect 42062 473618 42146 473854
rect 42382 473618 42414 473854
rect 41794 473534 42414 473618
rect 41794 473298 41826 473534
rect 42062 473298 42146 473534
rect 42382 473298 42414 473534
rect 77794 473618 77826 473854
rect 78062 473618 78146 473854
rect 78382 473618 78414 473854
rect 77794 473534 78414 473618
rect 77794 473298 77826 473534
rect 78062 473298 78146 473534
rect 78382 473298 78414 473534
rect 113794 473618 113826 473854
rect 114062 473618 114146 473854
rect 114382 473618 114414 473854
rect 113794 473534 114414 473618
rect 113794 473298 113826 473534
rect 114062 473298 114146 473534
rect 114382 473298 114414 473534
rect 149794 473618 149826 473854
rect 150062 473618 150146 473854
rect 150382 473618 150414 473854
rect 149794 473534 150414 473618
rect 149794 473298 149826 473534
rect 150062 473298 150146 473534
rect 150382 473298 150414 473534
rect 185794 473618 185826 473854
rect 186062 473618 186146 473854
rect 186382 473618 186414 473854
rect 185794 473534 186414 473618
rect 185794 473298 185826 473534
rect 186062 473298 186146 473534
rect 186382 473298 186414 473534
rect 221794 473618 221826 473854
rect 222062 473618 222146 473854
rect 222382 473618 222414 473854
rect 221794 473534 222414 473618
rect 221794 473298 221826 473534
rect 222062 473298 222146 473534
rect 222382 473298 222414 473534
rect 257794 473618 257826 473854
rect 258062 473618 258146 473854
rect 258382 473618 258414 473854
rect 257794 473534 258414 473618
rect 257794 473298 257826 473534
rect 258062 473298 258146 473534
rect 258382 473298 258414 473534
rect 293794 473618 293826 473854
rect 294062 473618 294146 473854
rect 294382 473618 294414 473854
rect 293794 473534 294414 473618
rect 293794 473298 293826 473534
rect 294062 473298 294146 473534
rect 294382 473298 294414 473534
rect 329794 473618 329826 473854
rect 330062 473618 330146 473854
rect 330382 473618 330414 473854
rect 329794 473534 330414 473618
rect 329794 473298 329826 473534
rect 330062 473298 330146 473534
rect 330382 473298 330414 473534
rect 365794 473618 365826 473854
rect 366062 473618 366146 473854
rect 366382 473618 366414 473854
rect 365794 473534 366414 473618
rect 365794 473298 365826 473534
rect 366062 473298 366146 473534
rect 366382 473298 366414 473534
rect 401794 473618 401826 473854
rect 402062 473618 402146 473854
rect 402382 473618 402414 473854
rect 401794 473534 402414 473618
rect 401794 473298 401826 473534
rect 402062 473298 402146 473534
rect 402382 473298 402414 473534
rect 437794 473618 437826 473854
rect 438062 473618 438146 473854
rect 438382 473618 438414 473854
rect 437794 473534 438414 473618
rect 437794 473298 437826 473534
rect 438062 473298 438146 473534
rect 438382 473298 438414 473534
rect 473794 473618 473826 473854
rect 474062 473618 474146 473854
rect 474382 473618 474414 473854
rect 473794 473534 474414 473618
rect 473794 473298 473826 473534
rect 474062 473298 474146 473534
rect 474382 473298 474414 473534
rect 509794 473618 509826 473854
rect 510062 473618 510146 473854
rect 510382 473618 510414 473854
rect 509794 473534 510414 473618
rect 509794 473298 509826 473534
rect 510062 473298 510146 473534
rect 510382 473298 510414 473534
rect 545794 473618 545826 473854
rect 546062 473618 546146 473854
rect 546382 473618 546414 473854
rect 545794 473534 546414 473618
rect 545794 473298 545826 473534
rect 546062 473298 546146 473534
rect 546382 473298 546414 473534
rect -2006 437854 -1386 473298
rect 582294 442354 582914 477798
rect 13166 442118 13198 442354
rect 13434 442118 13518 442354
rect 13754 442118 13786 442354
rect 13166 442034 13786 442118
rect 13166 441798 13198 442034
rect 13434 441798 13518 442034
rect 13754 441798 13786 442034
rect 167794 442118 167826 442354
rect 168062 442118 168146 442354
rect 168382 442118 168414 442354
rect 167794 442034 168414 442118
rect 167794 441798 167826 442034
rect 168062 441798 168146 442034
rect 168382 441798 168414 442034
rect 203794 442118 203826 442354
rect 204062 442118 204146 442354
rect 204382 442118 204414 442354
rect 203794 442034 204414 442118
rect 203794 441798 203826 442034
rect 204062 441798 204146 442034
rect 204382 441798 204414 442034
rect 239794 442118 239826 442354
rect 240062 442118 240146 442354
rect 240382 442118 240414 442354
rect 239794 442034 240414 442118
rect 239794 441798 239826 442034
rect 240062 441798 240146 442034
rect 240382 441798 240414 442034
rect 275794 442118 275826 442354
rect 276062 442118 276146 442354
rect 276382 442118 276414 442354
rect 275794 442034 276414 442118
rect 275794 441798 275826 442034
rect 276062 441798 276146 442034
rect 276382 441798 276414 442034
rect 311794 442118 311826 442354
rect 312062 442118 312146 442354
rect 312382 442118 312414 442354
rect 311794 442034 312414 442118
rect 311794 441798 311826 442034
rect 312062 441798 312146 442034
rect 312382 441798 312414 442034
rect 347794 442118 347826 442354
rect 348062 442118 348146 442354
rect 348382 442118 348414 442354
rect 347794 442034 348414 442118
rect 347794 441798 347826 442034
rect 348062 441798 348146 442034
rect 348382 441798 348414 442034
rect 383794 442118 383826 442354
rect 384062 442118 384146 442354
rect 384382 442118 384414 442354
rect 383794 442034 384414 442118
rect 383794 441798 383826 442034
rect 384062 441798 384146 442034
rect 384382 441798 384414 442034
rect 419794 442118 419826 442354
rect 420062 442118 420146 442354
rect 420382 442118 420414 442354
rect 419794 442034 420414 442118
rect 419794 441798 419826 442034
rect 420062 441798 420146 442034
rect 420382 441798 420414 442034
rect 563794 442118 563826 442354
rect 564062 442118 564146 442354
rect 564382 442118 564414 442354
rect 563794 442034 564414 442118
rect 563794 441798 563826 442034
rect 564062 441798 564146 442034
rect 564382 441798 564414 442034
rect 582294 442118 582326 442354
rect 582562 442118 582646 442354
rect 582882 442118 582914 442354
rect 582294 442034 582914 442118
rect 582294 441798 582326 442034
rect 582562 441798 582646 442034
rect 582882 441798 582914 442034
rect -2006 437618 -1974 437854
rect -1738 437618 -1654 437854
rect -1418 437618 -1386 437854
rect -2006 437534 -1386 437618
rect -2006 437298 -1974 437534
rect -1738 437298 -1654 437534
rect -1418 437298 -1386 437534
rect 5794 437618 5826 437854
rect 6062 437618 6146 437854
rect 6382 437618 6414 437854
rect 5794 437534 6414 437618
rect 5794 437298 5826 437534
rect 6062 437298 6146 437534
rect 6382 437298 6414 437534
rect 185794 437618 185826 437854
rect 186062 437618 186146 437854
rect 186382 437618 186414 437854
rect 185794 437534 186414 437618
rect 185794 437298 185826 437534
rect 186062 437298 186146 437534
rect 186382 437298 186414 437534
rect 221794 437618 221826 437854
rect 222062 437618 222146 437854
rect 222382 437618 222414 437854
rect 221794 437534 222414 437618
rect 221794 437298 221826 437534
rect 222062 437298 222146 437534
rect 222382 437298 222414 437534
rect 257794 437618 257826 437854
rect 258062 437618 258146 437854
rect 258382 437618 258414 437854
rect 257794 437534 258414 437618
rect 257794 437298 257826 437534
rect 258062 437298 258146 437534
rect 258382 437298 258414 437534
rect 293794 437618 293826 437854
rect 294062 437618 294146 437854
rect 294382 437618 294414 437854
rect 293794 437534 294414 437618
rect 293794 437298 293826 437534
rect 294062 437298 294146 437534
rect 294382 437298 294414 437534
rect 329794 437618 329826 437854
rect 330062 437618 330146 437854
rect 330382 437618 330414 437854
rect 329794 437534 330414 437618
rect 329794 437298 329826 437534
rect 330062 437298 330146 437534
rect 330382 437298 330414 437534
rect 365794 437618 365826 437854
rect 366062 437618 366146 437854
rect 366382 437618 366414 437854
rect 365794 437534 366414 437618
rect 365794 437298 365826 437534
rect 366062 437298 366146 437534
rect 366382 437298 366414 437534
rect 401794 437618 401826 437854
rect 402062 437618 402146 437854
rect 402382 437618 402414 437854
rect 401794 437534 402414 437618
rect 401794 437298 401826 437534
rect 402062 437298 402146 437534
rect 402382 437298 402414 437534
rect 570318 437618 570350 437854
rect 570586 437618 570670 437854
rect 570906 437618 570938 437854
rect 570318 437534 570938 437618
rect 570318 437298 570350 437534
rect 570586 437298 570670 437534
rect 570906 437298 570938 437534
rect -2006 401854 -1386 437298
rect 582294 406354 582914 441798
rect 13166 406118 13198 406354
rect 13434 406118 13518 406354
rect 13754 406118 13786 406354
rect 13166 406034 13786 406118
rect 13166 405798 13198 406034
rect 13434 405798 13518 406034
rect 13754 405798 13786 406034
rect 167794 406118 167826 406354
rect 168062 406118 168146 406354
rect 168382 406118 168414 406354
rect 167794 406034 168414 406118
rect 167794 405798 167826 406034
rect 168062 405798 168146 406034
rect 168382 405798 168414 406034
rect 203794 406118 203826 406354
rect 204062 406118 204146 406354
rect 204382 406118 204414 406354
rect 203794 406034 204414 406118
rect 203794 405798 203826 406034
rect 204062 405798 204146 406034
rect 204382 405798 204414 406034
rect 239794 406118 239826 406354
rect 240062 406118 240146 406354
rect 240382 406118 240414 406354
rect 239794 406034 240414 406118
rect 239794 405798 239826 406034
rect 240062 405798 240146 406034
rect 240382 405798 240414 406034
rect 275794 406118 275826 406354
rect 276062 406118 276146 406354
rect 276382 406118 276414 406354
rect 275794 406034 276414 406118
rect 275794 405798 275826 406034
rect 276062 405798 276146 406034
rect 276382 405798 276414 406034
rect 311794 406118 311826 406354
rect 312062 406118 312146 406354
rect 312382 406118 312414 406354
rect 311794 406034 312414 406118
rect 311794 405798 311826 406034
rect 312062 405798 312146 406034
rect 312382 405798 312414 406034
rect 347794 406118 347826 406354
rect 348062 406118 348146 406354
rect 348382 406118 348414 406354
rect 347794 406034 348414 406118
rect 347794 405798 347826 406034
rect 348062 405798 348146 406034
rect 348382 405798 348414 406034
rect 383794 406118 383826 406354
rect 384062 406118 384146 406354
rect 384382 406118 384414 406354
rect 383794 406034 384414 406118
rect 383794 405798 383826 406034
rect 384062 405798 384146 406034
rect 384382 405798 384414 406034
rect 419794 406118 419826 406354
rect 420062 406118 420146 406354
rect 420382 406118 420414 406354
rect 419794 406034 420414 406118
rect 419794 405798 419826 406034
rect 420062 405798 420146 406034
rect 420382 405798 420414 406034
rect 563794 406118 563826 406354
rect 564062 406118 564146 406354
rect 564382 406118 564414 406354
rect 563794 406034 564414 406118
rect 563794 405798 563826 406034
rect 564062 405798 564146 406034
rect 564382 405798 564414 406034
rect 582294 406118 582326 406354
rect 582562 406118 582646 406354
rect 582882 406118 582914 406354
rect 582294 406034 582914 406118
rect 582294 405798 582326 406034
rect 582562 405798 582646 406034
rect 582882 405798 582914 406034
rect -2006 401618 -1974 401854
rect -1738 401618 -1654 401854
rect -1418 401618 -1386 401854
rect -2006 401534 -1386 401618
rect -2006 401298 -1974 401534
rect -1738 401298 -1654 401534
rect -1418 401298 -1386 401534
rect 5794 401618 5826 401854
rect 6062 401618 6146 401854
rect 6382 401618 6414 401854
rect 5794 401534 6414 401618
rect 5794 401298 5826 401534
rect 6062 401298 6146 401534
rect 6382 401298 6414 401534
rect 185794 401618 185826 401854
rect 186062 401618 186146 401854
rect 186382 401618 186414 401854
rect 185794 401534 186414 401618
rect 185794 401298 185826 401534
rect 186062 401298 186146 401534
rect 186382 401298 186414 401534
rect 221794 401618 221826 401854
rect 222062 401618 222146 401854
rect 222382 401618 222414 401854
rect 221794 401534 222414 401618
rect 221794 401298 221826 401534
rect 222062 401298 222146 401534
rect 222382 401298 222414 401534
rect 257794 401618 257826 401854
rect 258062 401618 258146 401854
rect 258382 401618 258414 401854
rect 257794 401534 258414 401618
rect 257794 401298 257826 401534
rect 258062 401298 258146 401534
rect 258382 401298 258414 401534
rect 293794 401618 293826 401854
rect 294062 401618 294146 401854
rect 294382 401618 294414 401854
rect 293794 401534 294414 401618
rect 293794 401298 293826 401534
rect 294062 401298 294146 401534
rect 294382 401298 294414 401534
rect 329794 401618 329826 401854
rect 330062 401618 330146 401854
rect 330382 401618 330414 401854
rect 329794 401534 330414 401618
rect 329794 401298 329826 401534
rect 330062 401298 330146 401534
rect 330382 401298 330414 401534
rect 365794 401618 365826 401854
rect 366062 401618 366146 401854
rect 366382 401618 366414 401854
rect 365794 401534 366414 401618
rect 365794 401298 365826 401534
rect 366062 401298 366146 401534
rect 366382 401298 366414 401534
rect 401794 401618 401826 401854
rect 402062 401618 402146 401854
rect 402382 401618 402414 401854
rect 401794 401534 402414 401618
rect 401794 401298 401826 401534
rect 402062 401298 402146 401534
rect 402382 401298 402414 401534
rect 570318 401618 570350 401854
rect 570586 401618 570670 401854
rect 570906 401618 570938 401854
rect 570318 401534 570938 401618
rect 570318 401298 570350 401534
rect 570586 401298 570670 401534
rect 570906 401298 570938 401534
rect -2006 365854 -1386 401298
rect 582294 370354 582914 405798
rect 13166 370118 13198 370354
rect 13434 370118 13518 370354
rect 13754 370118 13786 370354
rect 13166 370034 13786 370118
rect 13166 369798 13198 370034
rect 13434 369798 13518 370034
rect 13754 369798 13786 370034
rect 167794 370118 167826 370354
rect 168062 370118 168146 370354
rect 168382 370118 168414 370354
rect 167794 370034 168414 370118
rect 167794 369798 167826 370034
rect 168062 369798 168146 370034
rect 168382 369798 168414 370034
rect 203794 370118 203826 370354
rect 204062 370118 204146 370354
rect 204382 370118 204414 370354
rect 203794 370034 204414 370118
rect 203794 369798 203826 370034
rect 204062 369798 204146 370034
rect 204382 369798 204414 370034
rect 239794 370118 239826 370354
rect 240062 370118 240146 370354
rect 240382 370118 240414 370354
rect 239794 370034 240414 370118
rect 239794 369798 239826 370034
rect 240062 369798 240146 370034
rect 240382 369798 240414 370034
rect 275794 370118 275826 370354
rect 276062 370118 276146 370354
rect 276382 370118 276414 370354
rect 275794 370034 276414 370118
rect 275794 369798 275826 370034
rect 276062 369798 276146 370034
rect 276382 369798 276414 370034
rect 311794 370118 311826 370354
rect 312062 370118 312146 370354
rect 312382 370118 312414 370354
rect 311794 370034 312414 370118
rect 311794 369798 311826 370034
rect 312062 369798 312146 370034
rect 312382 369798 312414 370034
rect 347794 370118 347826 370354
rect 348062 370118 348146 370354
rect 348382 370118 348414 370354
rect 347794 370034 348414 370118
rect 347794 369798 347826 370034
rect 348062 369798 348146 370034
rect 348382 369798 348414 370034
rect 383794 370118 383826 370354
rect 384062 370118 384146 370354
rect 384382 370118 384414 370354
rect 383794 370034 384414 370118
rect 383794 369798 383826 370034
rect 384062 369798 384146 370034
rect 384382 369798 384414 370034
rect 419794 370118 419826 370354
rect 420062 370118 420146 370354
rect 420382 370118 420414 370354
rect 419794 370034 420414 370118
rect 419794 369798 419826 370034
rect 420062 369798 420146 370034
rect 420382 369798 420414 370034
rect 563794 370118 563826 370354
rect 564062 370118 564146 370354
rect 564382 370118 564414 370354
rect 563794 370034 564414 370118
rect 563794 369798 563826 370034
rect 564062 369798 564146 370034
rect 564382 369798 564414 370034
rect 582294 370118 582326 370354
rect 582562 370118 582646 370354
rect 582882 370118 582914 370354
rect 582294 370034 582914 370118
rect 582294 369798 582326 370034
rect 582562 369798 582646 370034
rect 582882 369798 582914 370034
rect -2006 365618 -1974 365854
rect -1738 365618 -1654 365854
rect -1418 365618 -1386 365854
rect -2006 365534 -1386 365618
rect -2006 365298 -1974 365534
rect -1738 365298 -1654 365534
rect -1418 365298 -1386 365534
rect 5794 365618 5826 365854
rect 6062 365618 6146 365854
rect 6382 365618 6414 365854
rect 5794 365534 6414 365618
rect 5794 365298 5826 365534
rect 6062 365298 6146 365534
rect 6382 365298 6414 365534
rect 41794 365618 41826 365854
rect 42062 365618 42146 365854
rect 42382 365618 42414 365854
rect 41794 365534 42414 365618
rect 41794 365298 41826 365534
rect 42062 365298 42146 365534
rect 42382 365298 42414 365534
rect 77794 365618 77826 365854
rect 78062 365618 78146 365854
rect 78382 365618 78414 365854
rect 77794 365534 78414 365618
rect 77794 365298 77826 365534
rect 78062 365298 78146 365534
rect 78382 365298 78414 365534
rect 113794 365618 113826 365854
rect 114062 365618 114146 365854
rect 114382 365618 114414 365854
rect 113794 365534 114414 365618
rect 113794 365298 113826 365534
rect 114062 365298 114146 365534
rect 114382 365298 114414 365534
rect 149794 365618 149826 365854
rect 150062 365618 150146 365854
rect 150382 365618 150414 365854
rect 149794 365534 150414 365618
rect 149794 365298 149826 365534
rect 150062 365298 150146 365534
rect 150382 365298 150414 365534
rect 185794 365618 185826 365854
rect 186062 365618 186146 365854
rect 186382 365618 186414 365854
rect 185794 365534 186414 365618
rect 185794 365298 185826 365534
rect 186062 365298 186146 365534
rect 186382 365298 186414 365534
rect 221794 365618 221826 365854
rect 222062 365618 222146 365854
rect 222382 365618 222414 365854
rect 221794 365534 222414 365618
rect 221794 365298 221826 365534
rect 222062 365298 222146 365534
rect 222382 365298 222414 365534
rect 257794 365618 257826 365854
rect 258062 365618 258146 365854
rect 258382 365618 258414 365854
rect 257794 365534 258414 365618
rect 257794 365298 257826 365534
rect 258062 365298 258146 365534
rect 258382 365298 258414 365534
rect 293794 365618 293826 365854
rect 294062 365618 294146 365854
rect 294382 365618 294414 365854
rect 293794 365534 294414 365618
rect 293794 365298 293826 365534
rect 294062 365298 294146 365534
rect 294382 365298 294414 365534
rect 329794 365618 329826 365854
rect 330062 365618 330146 365854
rect 330382 365618 330414 365854
rect 329794 365534 330414 365618
rect 329794 365298 329826 365534
rect 330062 365298 330146 365534
rect 330382 365298 330414 365534
rect 365794 365618 365826 365854
rect 366062 365618 366146 365854
rect 366382 365618 366414 365854
rect 365794 365534 366414 365618
rect 365794 365298 365826 365534
rect 366062 365298 366146 365534
rect 366382 365298 366414 365534
rect 401794 365618 401826 365854
rect 402062 365618 402146 365854
rect 402382 365618 402414 365854
rect 401794 365534 402414 365618
rect 401794 365298 401826 365534
rect 402062 365298 402146 365534
rect 402382 365298 402414 365534
rect 437794 365618 437826 365854
rect 438062 365618 438146 365854
rect 438382 365618 438414 365854
rect 437794 365534 438414 365618
rect 437794 365298 437826 365534
rect 438062 365298 438146 365534
rect 438382 365298 438414 365534
rect 473794 365618 473826 365854
rect 474062 365618 474146 365854
rect 474382 365618 474414 365854
rect 473794 365534 474414 365618
rect 473794 365298 473826 365534
rect 474062 365298 474146 365534
rect 474382 365298 474414 365534
rect 509794 365618 509826 365854
rect 510062 365618 510146 365854
rect 510382 365618 510414 365854
rect 509794 365534 510414 365618
rect 509794 365298 509826 365534
rect 510062 365298 510146 365534
rect 510382 365298 510414 365534
rect 545794 365618 545826 365854
rect 546062 365618 546146 365854
rect 546382 365618 546414 365854
rect 545794 365534 546414 365618
rect 545794 365298 545826 365534
rect 546062 365298 546146 365534
rect 546382 365298 546414 365534
rect -2006 329854 -1386 365298
rect 582294 334354 582914 369798
rect 13166 334118 13198 334354
rect 13434 334118 13518 334354
rect 13754 334118 13786 334354
rect 13166 334034 13786 334118
rect 13166 333798 13198 334034
rect 13434 333798 13518 334034
rect 13754 333798 13786 334034
rect 167794 334118 167826 334354
rect 168062 334118 168146 334354
rect 168382 334118 168414 334354
rect 167794 334034 168414 334118
rect 167794 333798 167826 334034
rect 168062 333798 168146 334034
rect 168382 333798 168414 334034
rect 203794 334118 203826 334354
rect 204062 334118 204146 334354
rect 204382 334118 204414 334354
rect 203794 334034 204414 334118
rect 203794 333798 203826 334034
rect 204062 333798 204146 334034
rect 204382 333798 204414 334034
rect 239794 334118 239826 334354
rect 240062 334118 240146 334354
rect 240382 334118 240414 334354
rect 239794 334034 240414 334118
rect 239794 333798 239826 334034
rect 240062 333798 240146 334034
rect 240382 333798 240414 334034
rect 275794 334118 275826 334354
rect 276062 334118 276146 334354
rect 276382 334118 276414 334354
rect 275794 334034 276414 334118
rect 275794 333798 275826 334034
rect 276062 333798 276146 334034
rect 276382 333798 276414 334034
rect 311794 334118 311826 334354
rect 312062 334118 312146 334354
rect 312382 334118 312414 334354
rect 311794 334034 312414 334118
rect 311794 333798 311826 334034
rect 312062 333798 312146 334034
rect 312382 333798 312414 334034
rect 347794 334118 347826 334354
rect 348062 334118 348146 334354
rect 348382 334118 348414 334354
rect 347794 334034 348414 334118
rect 347794 333798 347826 334034
rect 348062 333798 348146 334034
rect 348382 333798 348414 334034
rect 383794 334118 383826 334354
rect 384062 334118 384146 334354
rect 384382 334118 384414 334354
rect 383794 334034 384414 334118
rect 383794 333798 383826 334034
rect 384062 333798 384146 334034
rect 384382 333798 384414 334034
rect 419794 334118 419826 334354
rect 420062 334118 420146 334354
rect 420382 334118 420414 334354
rect 419794 334034 420414 334118
rect 419794 333798 419826 334034
rect 420062 333798 420146 334034
rect 420382 333798 420414 334034
rect 563794 334118 563826 334354
rect 564062 334118 564146 334354
rect 564382 334118 564414 334354
rect 563794 334034 564414 334118
rect 563794 333798 563826 334034
rect 564062 333798 564146 334034
rect 564382 333798 564414 334034
rect 582294 334118 582326 334354
rect 582562 334118 582646 334354
rect 582882 334118 582914 334354
rect 582294 334034 582914 334118
rect 582294 333798 582326 334034
rect 582562 333798 582646 334034
rect 582882 333798 582914 334034
rect -2006 329618 -1974 329854
rect -1738 329618 -1654 329854
rect -1418 329618 -1386 329854
rect -2006 329534 -1386 329618
rect -2006 329298 -1974 329534
rect -1738 329298 -1654 329534
rect -1418 329298 -1386 329534
rect 5794 329618 5826 329854
rect 6062 329618 6146 329854
rect 6382 329618 6414 329854
rect 5794 329534 6414 329618
rect 5794 329298 5826 329534
rect 6062 329298 6146 329534
rect 6382 329298 6414 329534
rect 185794 329618 185826 329854
rect 186062 329618 186146 329854
rect 186382 329618 186414 329854
rect 185794 329534 186414 329618
rect 185794 329298 185826 329534
rect 186062 329298 186146 329534
rect 186382 329298 186414 329534
rect 221794 329618 221826 329854
rect 222062 329618 222146 329854
rect 222382 329618 222414 329854
rect 221794 329534 222414 329618
rect 221794 329298 221826 329534
rect 222062 329298 222146 329534
rect 222382 329298 222414 329534
rect 257794 329618 257826 329854
rect 258062 329618 258146 329854
rect 258382 329618 258414 329854
rect 257794 329534 258414 329618
rect 257794 329298 257826 329534
rect 258062 329298 258146 329534
rect 258382 329298 258414 329534
rect 293794 329618 293826 329854
rect 294062 329618 294146 329854
rect 294382 329618 294414 329854
rect 293794 329534 294414 329618
rect 293794 329298 293826 329534
rect 294062 329298 294146 329534
rect 294382 329298 294414 329534
rect 329794 329618 329826 329854
rect 330062 329618 330146 329854
rect 330382 329618 330414 329854
rect 329794 329534 330414 329618
rect 329794 329298 329826 329534
rect 330062 329298 330146 329534
rect 330382 329298 330414 329534
rect 365794 329618 365826 329854
rect 366062 329618 366146 329854
rect 366382 329618 366414 329854
rect 365794 329534 366414 329618
rect 365794 329298 365826 329534
rect 366062 329298 366146 329534
rect 366382 329298 366414 329534
rect 401794 329618 401826 329854
rect 402062 329618 402146 329854
rect 402382 329618 402414 329854
rect 401794 329534 402414 329618
rect 401794 329298 401826 329534
rect 402062 329298 402146 329534
rect 402382 329298 402414 329534
rect 570318 329618 570350 329854
rect 570586 329618 570670 329854
rect 570906 329618 570938 329854
rect 570318 329534 570938 329618
rect 570318 329298 570350 329534
rect 570586 329298 570670 329534
rect 570906 329298 570938 329534
rect -2006 293854 -1386 329298
rect 582294 298354 582914 333798
rect 13166 298118 13198 298354
rect 13434 298118 13518 298354
rect 13754 298118 13786 298354
rect 13166 298034 13786 298118
rect 13166 297798 13198 298034
rect 13434 297798 13518 298034
rect 13754 297798 13786 298034
rect 167794 298118 167826 298354
rect 168062 298118 168146 298354
rect 168382 298118 168414 298354
rect 167794 298034 168414 298118
rect 167794 297798 167826 298034
rect 168062 297798 168146 298034
rect 168382 297798 168414 298034
rect 203794 298118 203826 298354
rect 204062 298118 204146 298354
rect 204382 298118 204414 298354
rect 203794 298034 204414 298118
rect 203794 297798 203826 298034
rect 204062 297798 204146 298034
rect 204382 297798 204414 298034
rect 239794 298118 239826 298354
rect 240062 298118 240146 298354
rect 240382 298118 240414 298354
rect 239794 298034 240414 298118
rect 239794 297798 239826 298034
rect 240062 297798 240146 298034
rect 240382 297798 240414 298034
rect 275794 298118 275826 298354
rect 276062 298118 276146 298354
rect 276382 298118 276414 298354
rect 275794 298034 276414 298118
rect 275794 297798 275826 298034
rect 276062 297798 276146 298034
rect 276382 297798 276414 298034
rect 311794 298118 311826 298354
rect 312062 298118 312146 298354
rect 312382 298118 312414 298354
rect 311794 298034 312414 298118
rect 311794 297798 311826 298034
rect 312062 297798 312146 298034
rect 312382 297798 312414 298034
rect 347794 298118 347826 298354
rect 348062 298118 348146 298354
rect 348382 298118 348414 298354
rect 347794 298034 348414 298118
rect 347794 297798 347826 298034
rect 348062 297798 348146 298034
rect 348382 297798 348414 298034
rect 383794 298118 383826 298354
rect 384062 298118 384146 298354
rect 384382 298118 384414 298354
rect 383794 298034 384414 298118
rect 383794 297798 383826 298034
rect 384062 297798 384146 298034
rect 384382 297798 384414 298034
rect 419794 298118 419826 298354
rect 420062 298118 420146 298354
rect 420382 298118 420414 298354
rect 419794 298034 420414 298118
rect 419794 297798 419826 298034
rect 420062 297798 420146 298034
rect 420382 297798 420414 298034
rect 563794 298118 563826 298354
rect 564062 298118 564146 298354
rect 564382 298118 564414 298354
rect 563794 298034 564414 298118
rect 563794 297798 563826 298034
rect 564062 297798 564146 298034
rect 564382 297798 564414 298034
rect 582294 298118 582326 298354
rect 582562 298118 582646 298354
rect 582882 298118 582914 298354
rect 582294 298034 582914 298118
rect 582294 297798 582326 298034
rect 582562 297798 582646 298034
rect 582882 297798 582914 298034
rect -2006 293618 -1974 293854
rect -1738 293618 -1654 293854
rect -1418 293618 -1386 293854
rect -2006 293534 -1386 293618
rect -2006 293298 -1974 293534
rect -1738 293298 -1654 293534
rect -1418 293298 -1386 293534
rect 5794 293618 5826 293854
rect 6062 293618 6146 293854
rect 6382 293618 6414 293854
rect 5794 293534 6414 293618
rect 5794 293298 5826 293534
rect 6062 293298 6146 293534
rect 6382 293298 6414 293534
rect 185794 293618 185826 293854
rect 186062 293618 186146 293854
rect 186382 293618 186414 293854
rect 185794 293534 186414 293618
rect 185794 293298 185826 293534
rect 186062 293298 186146 293534
rect 186382 293298 186414 293534
rect 221794 293618 221826 293854
rect 222062 293618 222146 293854
rect 222382 293618 222414 293854
rect 221794 293534 222414 293618
rect 221794 293298 221826 293534
rect 222062 293298 222146 293534
rect 222382 293298 222414 293534
rect 257794 293618 257826 293854
rect 258062 293618 258146 293854
rect 258382 293618 258414 293854
rect 257794 293534 258414 293618
rect 257794 293298 257826 293534
rect 258062 293298 258146 293534
rect 258382 293298 258414 293534
rect 293794 293618 293826 293854
rect 294062 293618 294146 293854
rect 294382 293618 294414 293854
rect 293794 293534 294414 293618
rect 293794 293298 293826 293534
rect 294062 293298 294146 293534
rect 294382 293298 294414 293534
rect 329794 293618 329826 293854
rect 330062 293618 330146 293854
rect 330382 293618 330414 293854
rect 329794 293534 330414 293618
rect 329794 293298 329826 293534
rect 330062 293298 330146 293534
rect 330382 293298 330414 293534
rect 365794 293618 365826 293854
rect 366062 293618 366146 293854
rect 366382 293618 366414 293854
rect 365794 293534 366414 293618
rect 365794 293298 365826 293534
rect 366062 293298 366146 293534
rect 366382 293298 366414 293534
rect 401794 293618 401826 293854
rect 402062 293618 402146 293854
rect 402382 293618 402414 293854
rect 401794 293534 402414 293618
rect 401794 293298 401826 293534
rect 402062 293298 402146 293534
rect 402382 293298 402414 293534
rect 570318 293618 570350 293854
rect 570586 293618 570670 293854
rect 570906 293618 570938 293854
rect 570318 293534 570938 293618
rect 570318 293298 570350 293534
rect 570586 293298 570670 293534
rect 570906 293298 570938 293534
rect -2006 257854 -1386 293298
rect 582294 262354 582914 297798
rect 13166 262118 13198 262354
rect 13434 262118 13518 262354
rect 13754 262118 13786 262354
rect 13166 262034 13786 262118
rect 13166 261798 13198 262034
rect 13434 261798 13518 262034
rect 13754 261798 13786 262034
rect 167794 262118 167826 262354
rect 168062 262118 168146 262354
rect 168382 262118 168414 262354
rect 167794 262034 168414 262118
rect 167794 261798 167826 262034
rect 168062 261798 168146 262034
rect 168382 261798 168414 262034
rect 203794 262118 203826 262354
rect 204062 262118 204146 262354
rect 204382 262118 204414 262354
rect 203794 262034 204414 262118
rect 203794 261798 203826 262034
rect 204062 261798 204146 262034
rect 204382 261798 204414 262034
rect 239794 262118 239826 262354
rect 240062 262118 240146 262354
rect 240382 262118 240414 262354
rect 239794 262034 240414 262118
rect 239794 261798 239826 262034
rect 240062 261798 240146 262034
rect 240382 261798 240414 262034
rect 275794 262118 275826 262354
rect 276062 262118 276146 262354
rect 276382 262118 276414 262354
rect 275794 262034 276414 262118
rect 275794 261798 275826 262034
rect 276062 261798 276146 262034
rect 276382 261798 276414 262034
rect 311794 262118 311826 262354
rect 312062 262118 312146 262354
rect 312382 262118 312414 262354
rect 311794 262034 312414 262118
rect 311794 261798 311826 262034
rect 312062 261798 312146 262034
rect 312382 261798 312414 262034
rect 347794 262118 347826 262354
rect 348062 262118 348146 262354
rect 348382 262118 348414 262354
rect 347794 262034 348414 262118
rect 347794 261798 347826 262034
rect 348062 261798 348146 262034
rect 348382 261798 348414 262034
rect 383794 262118 383826 262354
rect 384062 262118 384146 262354
rect 384382 262118 384414 262354
rect 383794 262034 384414 262118
rect 383794 261798 383826 262034
rect 384062 261798 384146 262034
rect 384382 261798 384414 262034
rect 419794 262118 419826 262354
rect 420062 262118 420146 262354
rect 420382 262118 420414 262354
rect 419794 262034 420414 262118
rect 419794 261798 419826 262034
rect 420062 261798 420146 262034
rect 420382 261798 420414 262034
rect 563794 262118 563826 262354
rect 564062 262118 564146 262354
rect 564382 262118 564414 262354
rect 563794 262034 564414 262118
rect 563794 261798 563826 262034
rect 564062 261798 564146 262034
rect 564382 261798 564414 262034
rect 582294 262118 582326 262354
rect 582562 262118 582646 262354
rect 582882 262118 582914 262354
rect 582294 262034 582914 262118
rect 582294 261798 582326 262034
rect 582562 261798 582646 262034
rect 582882 261798 582914 262034
rect -2006 257618 -1974 257854
rect -1738 257618 -1654 257854
rect -1418 257618 -1386 257854
rect -2006 257534 -1386 257618
rect -2006 257298 -1974 257534
rect -1738 257298 -1654 257534
rect -1418 257298 -1386 257534
rect 5794 257618 5826 257854
rect 6062 257618 6146 257854
rect 6382 257618 6414 257854
rect 5794 257534 6414 257618
rect 5794 257298 5826 257534
rect 6062 257298 6146 257534
rect 6382 257298 6414 257534
rect 185794 257618 185826 257854
rect 186062 257618 186146 257854
rect 186382 257618 186414 257854
rect 185794 257534 186414 257618
rect 185794 257298 185826 257534
rect 186062 257298 186146 257534
rect 186382 257298 186414 257534
rect 221794 257618 221826 257854
rect 222062 257618 222146 257854
rect 222382 257618 222414 257854
rect 221794 257534 222414 257618
rect 221794 257298 221826 257534
rect 222062 257298 222146 257534
rect 222382 257298 222414 257534
rect 257794 257618 257826 257854
rect 258062 257618 258146 257854
rect 258382 257618 258414 257854
rect 257794 257534 258414 257618
rect 257794 257298 257826 257534
rect 258062 257298 258146 257534
rect 258382 257298 258414 257534
rect 293794 257618 293826 257854
rect 294062 257618 294146 257854
rect 294382 257618 294414 257854
rect 293794 257534 294414 257618
rect 293794 257298 293826 257534
rect 294062 257298 294146 257534
rect 294382 257298 294414 257534
rect 329794 257618 329826 257854
rect 330062 257618 330146 257854
rect 330382 257618 330414 257854
rect 329794 257534 330414 257618
rect 329794 257298 329826 257534
rect 330062 257298 330146 257534
rect 330382 257298 330414 257534
rect 365794 257618 365826 257854
rect 366062 257618 366146 257854
rect 366382 257618 366414 257854
rect 365794 257534 366414 257618
rect 365794 257298 365826 257534
rect 366062 257298 366146 257534
rect 366382 257298 366414 257534
rect 401794 257618 401826 257854
rect 402062 257618 402146 257854
rect 402382 257618 402414 257854
rect 401794 257534 402414 257618
rect 401794 257298 401826 257534
rect 402062 257298 402146 257534
rect 402382 257298 402414 257534
rect 570318 257618 570350 257854
rect 570586 257618 570670 257854
rect 570906 257618 570938 257854
rect 570318 257534 570938 257618
rect 570318 257298 570350 257534
rect 570586 257298 570670 257534
rect 570906 257298 570938 257534
rect -2006 221854 -1386 257298
rect 582294 226354 582914 261798
rect 23794 226118 23826 226354
rect 24062 226118 24146 226354
rect 24382 226118 24414 226354
rect 23794 226034 24414 226118
rect 23794 225798 23826 226034
rect 24062 225798 24146 226034
rect 24382 225798 24414 226034
rect 59794 226118 59826 226354
rect 60062 226118 60146 226354
rect 60382 226118 60414 226354
rect 59794 226034 60414 226118
rect 59794 225798 59826 226034
rect 60062 225798 60146 226034
rect 60382 225798 60414 226034
rect 95794 226118 95826 226354
rect 96062 226118 96146 226354
rect 96382 226118 96414 226354
rect 95794 226034 96414 226118
rect 95794 225798 95826 226034
rect 96062 225798 96146 226034
rect 96382 225798 96414 226034
rect 131794 226118 131826 226354
rect 132062 226118 132146 226354
rect 132382 226118 132414 226354
rect 131794 226034 132414 226118
rect 131794 225798 131826 226034
rect 132062 225798 132146 226034
rect 132382 225798 132414 226034
rect 167794 226118 167826 226354
rect 168062 226118 168146 226354
rect 168382 226118 168414 226354
rect 167794 226034 168414 226118
rect 167794 225798 167826 226034
rect 168062 225798 168146 226034
rect 168382 225798 168414 226034
rect 203794 226118 203826 226354
rect 204062 226118 204146 226354
rect 204382 226118 204414 226354
rect 203794 226034 204414 226118
rect 203794 225798 203826 226034
rect 204062 225798 204146 226034
rect 204382 225798 204414 226034
rect 239794 226118 239826 226354
rect 240062 226118 240146 226354
rect 240382 226118 240414 226354
rect 239794 226034 240414 226118
rect 239794 225798 239826 226034
rect 240062 225798 240146 226034
rect 240382 225798 240414 226034
rect 275794 226118 275826 226354
rect 276062 226118 276146 226354
rect 276382 226118 276414 226354
rect 275794 226034 276414 226118
rect 275794 225798 275826 226034
rect 276062 225798 276146 226034
rect 276382 225798 276414 226034
rect 311794 226118 311826 226354
rect 312062 226118 312146 226354
rect 312382 226118 312414 226354
rect 311794 226034 312414 226118
rect 311794 225798 311826 226034
rect 312062 225798 312146 226034
rect 312382 225798 312414 226034
rect 347794 226118 347826 226354
rect 348062 226118 348146 226354
rect 348382 226118 348414 226354
rect 347794 226034 348414 226118
rect 347794 225798 347826 226034
rect 348062 225798 348146 226034
rect 348382 225798 348414 226034
rect 383794 226118 383826 226354
rect 384062 226118 384146 226354
rect 384382 226118 384414 226354
rect 383794 226034 384414 226118
rect 383794 225798 383826 226034
rect 384062 225798 384146 226034
rect 384382 225798 384414 226034
rect 419794 226118 419826 226354
rect 420062 226118 420146 226354
rect 420382 226118 420414 226354
rect 419794 226034 420414 226118
rect 419794 225798 419826 226034
rect 420062 225798 420146 226034
rect 420382 225798 420414 226034
rect 455794 226118 455826 226354
rect 456062 226118 456146 226354
rect 456382 226118 456414 226354
rect 455794 226034 456414 226118
rect 455794 225798 455826 226034
rect 456062 225798 456146 226034
rect 456382 225798 456414 226034
rect 491794 226118 491826 226354
rect 492062 226118 492146 226354
rect 492382 226118 492414 226354
rect 491794 226034 492414 226118
rect 491794 225798 491826 226034
rect 492062 225798 492146 226034
rect 492382 225798 492414 226034
rect 527794 226118 527826 226354
rect 528062 226118 528146 226354
rect 528382 226118 528414 226354
rect 527794 226034 528414 226118
rect 527794 225798 527826 226034
rect 528062 225798 528146 226034
rect 528382 225798 528414 226034
rect 563794 226118 563826 226354
rect 564062 226118 564146 226354
rect 564382 226118 564414 226354
rect 563794 226034 564414 226118
rect 563794 225798 563826 226034
rect 564062 225798 564146 226034
rect 564382 225798 564414 226034
rect 582294 226118 582326 226354
rect 582562 226118 582646 226354
rect 582882 226118 582914 226354
rect 582294 226034 582914 226118
rect 582294 225798 582326 226034
rect 582562 225798 582646 226034
rect 582882 225798 582914 226034
rect -2006 221618 -1974 221854
rect -1738 221618 -1654 221854
rect -1418 221618 -1386 221854
rect -2006 221534 -1386 221618
rect -2006 221298 -1974 221534
rect -1738 221298 -1654 221534
rect -1418 221298 -1386 221534
rect 5794 221618 5826 221854
rect 6062 221618 6146 221854
rect 6382 221618 6414 221854
rect 5794 221534 6414 221618
rect 5794 221298 5826 221534
rect 6062 221298 6146 221534
rect 6382 221298 6414 221534
rect 185794 221618 185826 221854
rect 186062 221618 186146 221854
rect 186382 221618 186414 221854
rect 185794 221534 186414 221618
rect 185794 221298 185826 221534
rect 186062 221298 186146 221534
rect 186382 221298 186414 221534
rect 221794 221618 221826 221854
rect 222062 221618 222146 221854
rect 222382 221618 222414 221854
rect 221794 221534 222414 221618
rect 221794 221298 221826 221534
rect 222062 221298 222146 221534
rect 222382 221298 222414 221534
rect 257794 221618 257826 221854
rect 258062 221618 258146 221854
rect 258382 221618 258414 221854
rect 257794 221534 258414 221618
rect 257794 221298 257826 221534
rect 258062 221298 258146 221534
rect 258382 221298 258414 221534
rect 293794 221618 293826 221854
rect 294062 221618 294146 221854
rect 294382 221618 294414 221854
rect 293794 221534 294414 221618
rect 293794 221298 293826 221534
rect 294062 221298 294146 221534
rect 294382 221298 294414 221534
rect 329794 221618 329826 221854
rect 330062 221618 330146 221854
rect 330382 221618 330414 221854
rect 329794 221534 330414 221618
rect 329794 221298 329826 221534
rect 330062 221298 330146 221534
rect 330382 221298 330414 221534
rect 365794 221618 365826 221854
rect 366062 221618 366146 221854
rect 366382 221618 366414 221854
rect 365794 221534 366414 221618
rect 365794 221298 365826 221534
rect 366062 221298 366146 221534
rect 366382 221298 366414 221534
rect 401794 221618 401826 221854
rect 402062 221618 402146 221854
rect 402382 221618 402414 221854
rect 401794 221534 402414 221618
rect 401794 221298 401826 221534
rect 402062 221298 402146 221534
rect 402382 221298 402414 221534
rect 570318 221618 570350 221854
rect 570586 221618 570670 221854
rect 570906 221618 570938 221854
rect 570318 221534 570938 221618
rect 570318 221298 570350 221534
rect 570586 221298 570670 221534
rect 570906 221298 570938 221534
rect -2006 185854 -1386 221298
rect 582294 190354 582914 225798
rect 13166 190118 13198 190354
rect 13434 190118 13518 190354
rect 13754 190118 13786 190354
rect 13166 190034 13786 190118
rect 13166 189798 13198 190034
rect 13434 189798 13518 190034
rect 13754 189798 13786 190034
rect 167794 190118 167826 190354
rect 168062 190118 168146 190354
rect 168382 190118 168414 190354
rect 167794 190034 168414 190118
rect 167794 189798 167826 190034
rect 168062 189798 168146 190034
rect 168382 189798 168414 190034
rect 203794 190118 203826 190354
rect 204062 190118 204146 190354
rect 204382 190118 204414 190354
rect 203794 190034 204414 190118
rect 203794 189798 203826 190034
rect 204062 189798 204146 190034
rect 204382 189798 204414 190034
rect 239794 190118 239826 190354
rect 240062 190118 240146 190354
rect 240382 190118 240414 190354
rect 239794 190034 240414 190118
rect 239794 189798 239826 190034
rect 240062 189798 240146 190034
rect 240382 189798 240414 190034
rect 275794 190118 275826 190354
rect 276062 190118 276146 190354
rect 276382 190118 276414 190354
rect 275794 190034 276414 190118
rect 275794 189798 275826 190034
rect 276062 189798 276146 190034
rect 276382 189798 276414 190034
rect 311794 190118 311826 190354
rect 312062 190118 312146 190354
rect 312382 190118 312414 190354
rect 311794 190034 312414 190118
rect 311794 189798 311826 190034
rect 312062 189798 312146 190034
rect 312382 189798 312414 190034
rect 347794 190118 347826 190354
rect 348062 190118 348146 190354
rect 348382 190118 348414 190354
rect 347794 190034 348414 190118
rect 347794 189798 347826 190034
rect 348062 189798 348146 190034
rect 348382 189798 348414 190034
rect 383794 190118 383826 190354
rect 384062 190118 384146 190354
rect 384382 190118 384414 190354
rect 383794 190034 384414 190118
rect 383794 189798 383826 190034
rect 384062 189798 384146 190034
rect 384382 189798 384414 190034
rect 419794 190118 419826 190354
rect 420062 190118 420146 190354
rect 420382 190118 420414 190354
rect 419794 190034 420414 190118
rect 419794 189798 419826 190034
rect 420062 189798 420146 190034
rect 420382 189798 420414 190034
rect 563794 190118 563826 190354
rect 564062 190118 564146 190354
rect 564382 190118 564414 190354
rect 563794 190034 564414 190118
rect 563794 189798 563826 190034
rect 564062 189798 564146 190034
rect 564382 189798 564414 190034
rect 582294 190118 582326 190354
rect 582562 190118 582646 190354
rect 582882 190118 582914 190354
rect 582294 190034 582914 190118
rect 582294 189798 582326 190034
rect 582562 189798 582646 190034
rect 582882 189798 582914 190034
rect -2006 185618 -1974 185854
rect -1738 185618 -1654 185854
rect -1418 185618 -1386 185854
rect -2006 185534 -1386 185618
rect -2006 185298 -1974 185534
rect -1738 185298 -1654 185534
rect -1418 185298 -1386 185534
rect 5794 185618 5826 185854
rect 6062 185618 6146 185854
rect 6382 185618 6414 185854
rect 5794 185534 6414 185618
rect 5794 185298 5826 185534
rect 6062 185298 6146 185534
rect 6382 185298 6414 185534
rect 185794 185618 185826 185854
rect 186062 185618 186146 185854
rect 186382 185618 186414 185854
rect 185794 185534 186414 185618
rect 185794 185298 185826 185534
rect 186062 185298 186146 185534
rect 186382 185298 186414 185534
rect 221794 185618 221826 185854
rect 222062 185618 222146 185854
rect 222382 185618 222414 185854
rect 221794 185534 222414 185618
rect 221794 185298 221826 185534
rect 222062 185298 222146 185534
rect 222382 185298 222414 185534
rect 257794 185618 257826 185854
rect 258062 185618 258146 185854
rect 258382 185618 258414 185854
rect 257794 185534 258414 185618
rect 257794 185298 257826 185534
rect 258062 185298 258146 185534
rect 258382 185298 258414 185534
rect 293794 185618 293826 185854
rect 294062 185618 294146 185854
rect 294382 185618 294414 185854
rect 293794 185534 294414 185618
rect 293794 185298 293826 185534
rect 294062 185298 294146 185534
rect 294382 185298 294414 185534
rect 329794 185618 329826 185854
rect 330062 185618 330146 185854
rect 330382 185618 330414 185854
rect 329794 185534 330414 185618
rect 329794 185298 329826 185534
rect 330062 185298 330146 185534
rect 330382 185298 330414 185534
rect 365794 185618 365826 185854
rect 366062 185618 366146 185854
rect 366382 185618 366414 185854
rect 365794 185534 366414 185618
rect 365794 185298 365826 185534
rect 366062 185298 366146 185534
rect 366382 185298 366414 185534
rect 401794 185618 401826 185854
rect 402062 185618 402146 185854
rect 402382 185618 402414 185854
rect 401794 185534 402414 185618
rect 401794 185298 401826 185534
rect 402062 185298 402146 185534
rect 402382 185298 402414 185534
rect 570318 185618 570350 185854
rect 570586 185618 570670 185854
rect 570906 185618 570938 185854
rect 570318 185534 570938 185618
rect 570318 185298 570350 185534
rect 570586 185298 570670 185534
rect 570906 185298 570938 185534
rect -2006 149854 -1386 185298
rect 582294 154354 582914 189798
rect 13166 154118 13198 154354
rect 13434 154118 13518 154354
rect 13754 154118 13786 154354
rect 13166 154034 13786 154118
rect 13166 153798 13198 154034
rect 13434 153798 13518 154034
rect 13754 153798 13786 154034
rect 167794 154118 167826 154354
rect 168062 154118 168146 154354
rect 168382 154118 168414 154354
rect 167794 154034 168414 154118
rect 167794 153798 167826 154034
rect 168062 153798 168146 154034
rect 168382 153798 168414 154034
rect 203794 154118 203826 154354
rect 204062 154118 204146 154354
rect 204382 154118 204414 154354
rect 203794 154034 204414 154118
rect 203794 153798 203826 154034
rect 204062 153798 204146 154034
rect 204382 153798 204414 154034
rect 239794 154118 239826 154354
rect 240062 154118 240146 154354
rect 240382 154118 240414 154354
rect 239794 154034 240414 154118
rect 239794 153798 239826 154034
rect 240062 153798 240146 154034
rect 240382 153798 240414 154034
rect 275794 154118 275826 154354
rect 276062 154118 276146 154354
rect 276382 154118 276414 154354
rect 275794 154034 276414 154118
rect 275794 153798 275826 154034
rect 276062 153798 276146 154034
rect 276382 153798 276414 154034
rect 311794 154118 311826 154354
rect 312062 154118 312146 154354
rect 312382 154118 312414 154354
rect 311794 154034 312414 154118
rect 311794 153798 311826 154034
rect 312062 153798 312146 154034
rect 312382 153798 312414 154034
rect 347794 154118 347826 154354
rect 348062 154118 348146 154354
rect 348382 154118 348414 154354
rect 347794 154034 348414 154118
rect 347794 153798 347826 154034
rect 348062 153798 348146 154034
rect 348382 153798 348414 154034
rect 383794 154118 383826 154354
rect 384062 154118 384146 154354
rect 384382 154118 384414 154354
rect 383794 154034 384414 154118
rect 383794 153798 383826 154034
rect 384062 153798 384146 154034
rect 384382 153798 384414 154034
rect 419794 154118 419826 154354
rect 420062 154118 420146 154354
rect 420382 154118 420414 154354
rect 419794 154034 420414 154118
rect 419794 153798 419826 154034
rect 420062 153798 420146 154034
rect 420382 153798 420414 154034
rect 563794 154118 563826 154354
rect 564062 154118 564146 154354
rect 564382 154118 564414 154354
rect 563794 154034 564414 154118
rect 563794 153798 563826 154034
rect 564062 153798 564146 154034
rect 564382 153798 564414 154034
rect 582294 154118 582326 154354
rect 582562 154118 582646 154354
rect 582882 154118 582914 154354
rect 582294 154034 582914 154118
rect 582294 153798 582326 154034
rect 582562 153798 582646 154034
rect 582882 153798 582914 154034
rect -2006 149618 -1974 149854
rect -1738 149618 -1654 149854
rect -1418 149618 -1386 149854
rect -2006 149534 -1386 149618
rect -2006 149298 -1974 149534
rect -1738 149298 -1654 149534
rect -1418 149298 -1386 149534
rect 5794 149618 5826 149854
rect 6062 149618 6146 149854
rect 6382 149618 6414 149854
rect 5794 149534 6414 149618
rect 5794 149298 5826 149534
rect 6062 149298 6146 149534
rect 6382 149298 6414 149534
rect 185794 149618 185826 149854
rect 186062 149618 186146 149854
rect 186382 149618 186414 149854
rect 185794 149534 186414 149618
rect 185794 149298 185826 149534
rect 186062 149298 186146 149534
rect 186382 149298 186414 149534
rect 221794 149618 221826 149854
rect 222062 149618 222146 149854
rect 222382 149618 222414 149854
rect 221794 149534 222414 149618
rect 221794 149298 221826 149534
rect 222062 149298 222146 149534
rect 222382 149298 222414 149534
rect 257794 149618 257826 149854
rect 258062 149618 258146 149854
rect 258382 149618 258414 149854
rect 257794 149534 258414 149618
rect 257794 149298 257826 149534
rect 258062 149298 258146 149534
rect 258382 149298 258414 149534
rect 293794 149618 293826 149854
rect 294062 149618 294146 149854
rect 294382 149618 294414 149854
rect 293794 149534 294414 149618
rect 293794 149298 293826 149534
rect 294062 149298 294146 149534
rect 294382 149298 294414 149534
rect 329794 149618 329826 149854
rect 330062 149618 330146 149854
rect 330382 149618 330414 149854
rect 329794 149534 330414 149618
rect 329794 149298 329826 149534
rect 330062 149298 330146 149534
rect 330382 149298 330414 149534
rect 365794 149618 365826 149854
rect 366062 149618 366146 149854
rect 366382 149618 366414 149854
rect 365794 149534 366414 149618
rect 365794 149298 365826 149534
rect 366062 149298 366146 149534
rect 366382 149298 366414 149534
rect 401794 149618 401826 149854
rect 402062 149618 402146 149854
rect 402382 149618 402414 149854
rect 401794 149534 402414 149618
rect 401794 149298 401826 149534
rect 402062 149298 402146 149534
rect 402382 149298 402414 149534
rect 570318 149618 570350 149854
rect 570586 149618 570670 149854
rect 570906 149618 570938 149854
rect 570318 149534 570938 149618
rect 570318 149298 570350 149534
rect 570586 149298 570670 149534
rect 570906 149298 570938 149534
rect -2006 113854 -1386 149298
rect 582294 118354 582914 153798
rect 23794 118118 23826 118354
rect 24062 118118 24146 118354
rect 24382 118118 24414 118354
rect 23794 118034 24414 118118
rect 23794 117798 23826 118034
rect 24062 117798 24146 118034
rect 24382 117798 24414 118034
rect 59794 118118 59826 118354
rect 60062 118118 60146 118354
rect 60382 118118 60414 118354
rect 59794 118034 60414 118118
rect 59794 117798 59826 118034
rect 60062 117798 60146 118034
rect 60382 117798 60414 118034
rect 95794 118118 95826 118354
rect 96062 118118 96146 118354
rect 96382 118118 96414 118354
rect 95794 118034 96414 118118
rect 95794 117798 95826 118034
rect 96062 117798 96146 118034
rect 96382 117798 96414 118034
rect 131794 118118 131826 118354
rect 132062 118118 132146 118354
rect 132382 118118 132414 118354
rect 131794 118034 132414 118118
rect 131794 117798 131826 118034
rect 132062 117798 132146 118034
rect 132382 117798 132414 118034
rect 167794 118118 167826 118354
rect 168062 118118 168146 118354
rect 168382 118118 168414 118354
rect 167794 118034 168414 118118
rect 167794 117798 167826 118034
rect 168062 117798 168146 118034
rect 168382 117798 168414 118034
rect 203794 118118 203826 118354
rect 204062 118118 204146 118354
rect 204382 118118 204414 118354
rect 203794 118034 204414 118118
rect 203794 117798 203826 118034
rect 204062 117798 204146 118034
rect 204382 117798 204414 118034
rect 239794 118118 239826 118354
rect 240062 118118 240146 118354
rect 240382 118118 240414 118354
rect 239794 118034 240414 118118
rect 239794 117798 239826 118034
rect 240062 117798 240146 118034
rect 240382 117798 240414 118034
rect 275794 118118 275826 118354
rect 276062 118118 276146 118354
rect 276382 118118 276414 118354
rect 275794 118034 276414 118118
rect 275794 117798 275826 118034
rect 276062 117798 276146 118034
rect 276382 117798 276414 118034
rect 311794 118118 311826 118354
rect 312062 118118 312146 118354
rect 312382 118118 312414 118354
rect 311794 118034 312414 118118
rect 311794 117798 311826 118034
rect 312062 117798 312146 118034
rect 312382 117798 312414 118034
rect 347794 118118 347826 118354
rect 348062 118118 348146 118354
rect 348382 118118 348414 118354
rect 347794 118034 348414 118118
rect 347794 117798 347826 118034
rect 348062 117798 348146 118034
rect 348382 117798 348414 118034
rect 383794 118118 383826 118354
rect 384062 118118 384146 118354
rect 384382 118118 384414 118354
rect 383794 118034 384414 118118
rect 383794 117798 383826 118034
rect 384062 117798 384146 118034
rect 384382 117798 384414 118034
rect 419794 118118 419826 118354
rect 420062 118118 420146 118354
rect 420382 118118 420414 118354
rect 419794 118034 420414 118118
rect 419794 117798 419826 118034
rect 420062 117798 420146 118034
rect 420382 117798 420414 118034
rect 455794 118118 455826 118354
rect 456062 118118 456146 118354
rect 456382 118118 456414 118354
rect 455794 118034 456414 118118
rect 455794 117798 455826 118034
rect 456062 117798 456146 118034
rect 456382 117798 456414 118034
rect 491794 118118 491826 118354
rect 492062 118118 492146 118354
rect 492382 118118 492414 118354
rect 491794 118034 492414 118118
rect 491794 117798 491826 118034
rect 492062 117798 492146 118034
rect 492382 117798 492414 118034
rect 527794 118118 527826 118354
rect 528062 118118 528146 118354
rect 528382 118118 528414 118354
rect 527794 118034 528414 118118
rect 527794 117798 527826 118034
rect 528062 117798 528146 118034
rect 528382 117798 528414 118034
rect 563794 118118 563826 118354
rect 564062 118118 564146 118354
rect 564382 118118 564414 118354
rect 563794 118034 564414 118118
rect 563794 117798 563826 118034
rect 564062 117798 564146 118034
rect 564382 117798 564414 118034
rect 582294 118118 582326 118354
rect 582562 118118 582646 118354
rect 582882 118118 582914 118354
rect 582294 118034 582914 118118
rect 582294 117798 582326 118034
rect 582562 117798 582646 118034
rect 582882 117798 582914 118034
rect -2006 113618 -1974 113854
rect -1738 113618 -1654 113854
rect -1418 113618 -1386 113854
rect -2006 113534 -1386 113618
rect -2006 113298 -1974 113534
rect -1738 113298 -1654 113534
rect -1418 113298 -1386 113534
rect 5794 113618 5826 113854
rect 6062 113618 6146 113854
rect 6382 113618 6414 113854
rect 5794 113534 6414 113618
rect 5794 113298 5826 113534
rect 6062 113298 6146 113534
rect 6382 113298 6414 113534
rect 41794 113715 42414 113886
rect 41794 113479 41826 113715
rect 42062 113479 42146 113715
rect 42382 113479 42414 113715
rect 41794 113308 42414 113479
rect 77794 113715 78414 113886
rect 77794 113479 77826 113715
rect 78062 113479 78146 113715
rect 78382 113479 78414 113715
rect 77794 113308 78414 113479
rect 113794 113715 114414 113886
rect 113794 113479 113826 113715
rect 114062 113479 114146 113715
rect 114382 113479 114414 113715
rect 113794 113308 114414 113479
rect 149794 113715 150414 113886
rect 149794 113479 149826 113715
rect 150062 113479 150146 113715
rect 150382 113479 150414 113715
rect 149794 113308 150414 113479
rect 293794 113618 293826 113854
rect 294062 113618 294146 113854
rect 294382 113618 294414 113854
rect 293794 113534 294414 113618
rect 293794 113298 293826 113534
rect 294062 113298 294146 113534
rect 294382 113298 294414 113534
rect 401794 113618 401826 113854
rect 402062 113618 402146 113854
rect 402382 113618 402414 113854
rect 401794 113534 402414 113618
rect 401794 113298 401826 113534
rect 402062 113298 402146 113534
rect 402382 113298 402414 113534
rect 437794 113715 438414 113886
rect 437794 113479 437826 113715
rect 438062 113479 438146 113715
rect 438382 113479 438414 113715
rect 437794 113308 438414 113479
rect 473794 113715 474414 113886
rect 473794 113479 473826 113715
rect 474062 113479 474146 113715
rect 474382 113479 474414 113715
rect 473794 113308 474414 113479
rect 509794 113715 510414 113886
rect 509794 113479 509826 113715
rect 510062 113479 510146 113715
rect 510382 113479 510414 113715
rect 509794 113308 510414 113479
rect 545794 113715 546414 113886
rect 545794 113479 545826 113715
rect 546062 113479 546146 113715
rect 546382 113479 546414 113715
rect 545794 113308 546414 113479
rect -2006 77854 -1386 113298
rect 582294 82354 582914 117798
rect 13166 82118 13198 82354
rect 13434 82118 13518 82354
rect 13754 82118 13786 82354
rect 13166 82034 13786 82118
rect 13166 81798 13198 82034
rect 13434 81798 13518 82034
rect 13754 81798 13786 82034
rect 167794 82118 167826 82354
rect 168062 82118 168146 82354
rect 168382 82118 168414 82354
rect 167794 82034 168414 82118
rect 167794 81798 167826 82034
rect 168062 81798 168146 82034
rect 168382 81798 168414 82034
rect 291558 82118 291590 82354
rect 291826 82118 291910 82354
rect 292146 82118 292178 82354
rect 291558 82034 292178 82118
rect 291558 81798 291590 82034
rect 291826 81798 291910 82034
rect 292146 81798 292178 82034
rect 419794 82118 419826 82354
rect 420062 82118 420146 82354
rect 420382 82118 420414 82354
rect 419794 82034 420414 82118
rect 419794 81798 419826 82034
rect 420062 81798 420146 82034
rect 420382 81798 420414 82034
rect 563794 82118 563826 82354
rect 564062 82118 564146 82354
rect 564382 82118 564414 82354
rect 563794 82034 564414 82118
rect 563794 81798 563826 82034
rect 564062 81798 564146 82034
rect 564382 81798 564414 82034
rect 582294 82118 582326 82354
rect 582562 82118 582646 82354
rect 582882 82118 582914 82354
rect 582294 82034 582914 82118
rect 582294 81798 582326 82034
rect 582562 81798 582646 82034
rect 582882 81798 582914 82034
rect -2006 77618 -1974 77854
rect -1738 77618 -1654 77854
rect -1418 77618 -1386 77854
rect -2006 77534 -1386 77618
rect -2006 77298 -1974 77534
rect -1738 77298 -1654 77534
rect -1418 77298 -1386 77534
rect 5794 77618 5826 77854
rect 6062 77618 6146 77854
rect 6382 77618 6414 77854
rect 5794 77534 6414 77618
rect 5794 77298 5826 77534
rect 6062 77298 6146 77534
rect 6382 77298 6414 77534
rect 173062 77618 173094 77854
rect 173330 77618 173414 77854
rect 173650 77618 173682 77854
rect 173062 77534 173682 77618
rect 173062 77298 173094 77534
rect 173330 77298 173414 77534
rect 173650 77298 173682 77534
rect 293794 77618 293826 77854
rect 294062 77618 294146 77854
rect 294382 77618 294414 77854
rect 293794 77534 294414 77618
rect 293794 77298 293826 77534
rect 294062 77298 294146 77534
rect 294382 77298 294414 77534
rect 401794 77618 401826 77854
rect 402062 77618 402146 77854
rect 402382 77618 402414 77854
rect 401794 77534 402414 77618
rect 401794 77298 401826 77534
rect 402062 77298 402146 77534
rect 402382 77298 402414 77534
rect 570318 77618 570350 77854
rect 570586 77618 570670 77854
rect 570906 77618 570938 77854
rect 570318 77534 570938 77618
rect 570318 77298 570350 77534
rect 570586 77298 570670 77534
rect 570906 77298 570938 77534
rect -2006 41854 -1386 77298
rect 582294 46354 582914 81798
rect 13166 46118 13198 46354
rect 13434 46118 13518 46354
rect 13754 46118 13786 46354
rect 13166 46034 13786 46118
rect 13166 45798 13198 46034
rect 13434 45798 13518 46034
rect 13754 45798 13786 46034
rect 167794 46118 167826 46354
rect 168062 46118 168146 46354
rect 168382 46118 168414 46354
rect 167794 46034 168414 46118
rect 167794 45798 167826 46034
rect 168062 45798 168146 46034
rect 168382 45798 168414 46034
rect 291558 46118 291590 46354
rect 291826 46118 291910 46354
rect 292146 46118 292178 46354
rect 291558 46034 292178 46118
rect 291558 45798 291590 46034
rect 291826 45798 291910 46034
rect 292146 45798 292178 46034
rect 419794 46118 419826 46354
rect 420062 46118 420146 46354
rect 420382 46118 420414 46354
rect 419794 46034 420414 46118
rect 419794 45798 419826 46034
rect 420062 45798 420146 46034
rect 420382 45798 420414 46034
rect 563794 46118 563826 46354
rect 564062 46118 564146 46354
rect 564382 46118 564414 46354
rect 563794 46034 564414 46118
rect 563794 45798 563826 46034
rect 564062 45798 564146 46034
rect 564382 45798 564414 46034
rect 582294 46118 582326 46354
rect 582562 46118 582646 46354
rect 582882 46118 582914 46354
rect 582294 46034 582914 46118
rect 582294 45798 582326 46034
rect 582562 45798 582646 46034
rect 582882 45798 582914 46034
rect -2006 41618 -1974 41854
rect -1738 41618 -1654 41854
rect -1418 41618 -1386 41854
rect -2006 41534 -1386 41618
rect -2006 41298 -1974 41534
rect -1738 41298 -1654 41534
rect -1418 41298 -1386 41534
rect 5794 41618 5826 41854
rect 6062 41618 6146 41854
rect 6382 41618 6414 41854
rect 5794 41534 6414 41618
rect 5794 41298 5826 41534
rect 6062 41298 6146 41534
rect 6382 41298 6414 41534
rect 173062 41618 173094 41854
rect 173330 41618 173414 41854
rect 173650 41618 173682 41854
rect 173062 41534 173682 41618
rect 173062 41298 173094 41534
rect 173330 41298 173414 41534
rect 173650 41298 173682 41534
rect 293794 41618 293826 41854
rect 294062 41618 294146 41854
rect 294382 41618 294414 41854
rect 293794 41534 294414 41618
rect 293794 41298 293826 41534
rect 294062 41298 294146 41534
rect 294382 41298 294414 41534
rect 401794 41618 401826 41854
rect 402062 41618 402146 41854
rect 402382 41618 402414 41854
rect 401794 41534 402414 41618
rect 401794 41298 401826 41534
rect 402062 41298 402146 41534
rect 402382 41298 402414 41534
rect 570318 41618 570350 41854
rect 570586 41618 570670 41854
rect 570906 41618 570938 41854
rect 570318 41534 570938 41618
rect 570318 41298 570350 41534
rect 570586 41298 570670 41534
rect 570906 41298 570938 41534
rect -2006 5854 -1386 41298
rect 582294 10354 582914 45798
rect 23794 10118 23826 10354
rect 24062 10118 24146 10354
rect 24382 10118 24414 10354
rect 23794 10034 24414 10118
rect 23794 9798 23826 10034
rect 24062 9798 24146 10034
rect 24382 9798 24414 10034
rect 59794 10118 59826 10354
rect 60062 10118 60146 10354
rect 60382 10118 60414 10354
rect 59794 10034 60414 10118
rect 59794 9798 59826 10034
rect 60062 9798 60146 10034
rect 60382 9798 60414 10034
rect 95794 10118 95826 10354
rect 96062 10118 96146 10354
rect 96382 10118 96414 10354
rect 95794 10034 96414 10118
rect 95794 9798 95826 10034
rect 96062 9798 96146 10034
rect 96382 9798 96414 10034
rect 131794 10118 131826 10354
rect 132062 10118 132146 10354
rect 132382 10118 132414 10354
rect 131794 10034 132414 10118
rect 131794 9798 131826 10034
rect 132062 9798 132146 10034
rect 132382 9798 132414 10034
rect 167794 10118 167826 10354
rect 168062 10118 168146 10354
rect 168382 10118 168414 10354
rect 167794 10034 168414 10118
rect 167794 9798 167826 10034
rect 168062 9798 168146 10034
rect 168382 9798 168414 10034
rect 203794 10118 203826 10354
rect 204062 10118 204146 10354
rect 204382 10118 204414 10354
rect 203794 10034 204414 10118
rect 203794 9798 203826 10034
rect 204062 9798 204146 10034
rect 204382 9798 204414 10034
rect 239794 10118 239826 10354
rect 240062 10118 240146 10354
rect 240382 10118 240414 10354
rect 239794 10034 240414 10118
rect 239794 9798 239826 10034
rect 240062 9798 240146 10034
rect 240382 9798 240414 10034
rect 275794 10118 275826 10354
rect 276062 10118 276146 10354
rect 276382 10118 276414 10354
rect 275794 10034 276414 10118
rect 275794 9798 275826 10034
rect 276062 9798 276146 10034
rect 276382 9798 276414 10034
rect 311794 10118 311826 10354
rect 312062 10118 312146 10354
rect 312382 10118 312414 10354
rect 311794 10034 312414 10118
rect 311794 9798 311826 10034
rect 312062 9798 312146 10034
rect 312382 9798 312414 10034
rect 347794 10118 347826 10354
rect 348062 10118 348146 10354
rect 348382 10118 348414 10354
rect 347794 10034 348414 10118
rect 347794 9798 347826 10034
rect 348062 9798 348146 10034
rect 348382 9798 348414 10034
rect 383794 10118 383826 10354
rect 384062 10118 384146 10354
rect 384382 10118 384414 10354
rect 383794 10034 384414 10118
rect 383794 9798 383826 10034
rect 384062 9798 384146 10034
rect 384382 9798 384414 10034
rect 419794 10118 419826 10354
rect 420062 10118 420146 10354
rect 420382 10118 420414 10354
rect 419794 10034 420414 10118
rect 419794 9798 419826 10034
rect 420062 9798 420146 10034
rect 420382 9798 420414 10034
rect 455794 10118 455826 10354
rect 456062 10118 456146 10354
rect 456382 10118 456414 10354
rect 455794 10034 456414 10118
rect 455794 9798 455826 10034
rect 456062 9798 456146 10034
rect 456382 9798 456414 10034
rect 491794 10118 491826 10354
rect 492062 10118 492146 10354
rect 492382 10118 492414 10354
rect 491794 10034 492414 10118
rect 491794 9798 491826 10034
rect 492062 9798 492146 10034
rect 492382 9798 492414 10034
rect 527794 10118 527826 10354
rect 528062 10118 528146 10354
rect 528382 10118 528414 10354
rect 527794 10034 528414 10118
rect 527794 9798 527826 10034
rect 528062 9798 528146 10034
rect 528382 9798 528414 10034
rect 563794 10118 563826 10354
rect 564062 10118 564146 10354
rect 564382 10118 564414 10354
rect 563794 10034 564414 10118
rect 563794 9798 563826 10034
rect 564062 9798 564146 10034
rect 564382 9798 564414 10034
rect 582294 10118 582326 10354
rect 582562 10118 582646 10354
rect 582882 10118 582914 10354
rect 582294 10034 582914 10118
rect 582294 9798 582326 10034
rect 582562 9798 582646 10034
rect 582882 9798 582914 10034
rect -2006 5618 -1974 5854
rect -1738 5618 -1654 5854
rect -1418 5618 -1386 5854
rect -2006 5534 -1386 5618
rect -2006 5298 -1974 5534
rect -1738 5298 -1654 5534
rect -1418 5298 -1386 5534
rect -2006 -346 -1386 5298
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect 582294 -1306 582914 9798
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 689854 585930 704282
rect 585310 689618 585342 689854
rect 585578 689618 585662 689854
rect 585898 689618 585930 689854
rect 585310 689534 585930 689618
rect 585310 689298 585342 689534
rect 585578 689298 585662 689534
rect 585898 689298 585930 689534
rect 585310 653854 585930 689298
rect 585310 653618 585342 653854
rect 585578 653618 585662 653854
rect 585898 653618 585930 653854
rect 585310 653534 585930 653618
rect 585310 653298 585342 653534
rect 585578 653298 585662 653534
rect 585898 653298 585930 653534
rect 585310 617854 585930 653298
rect 585310 617618 585342 617854
rect 585578 617618 585662 617854
rect 585898 617618 585930 617854
rect 585310 617534 585930 617618
rect 585310 617298 585342 617534
rect 585578 617298 585662 617534
rect 585898 617298 585930 617534
rect 585310 581854 585930 617298
rect 585310 581618 585342 581854
rect 585578 581618 585662 581854
rect 585898 581618 585930 581854
rect 585310 581534 585930 581618
rect 585310 581298 585342 581534
rect 585578 581298 585662 581534
rect 585898 581298 585930 581534
rect 585310 545854 585930 581298
rect 585310 545618 585342 545854
rect 585578 545618 585662 545854
rect 585898 545618 585930 545854
rect 585310 545534 585930 545618
rect 585310 545298 585342 545534
rect 585578 545298 585662 545534
rect 585898 545298 585930 545534
rect 585310 509854 585930 545298
rect 585310 509618 585342 509854
rect 585578 509618 585662 509854
rect 585898 509618 585930 509854
rect 585310 509534 585930 509618
rect 585310 509298 585342 509534
rect 585578 509298 585662 509534
rect 585898 509298 585930 509534
rect 585310 473854 585930 509298
rect 585310 473618 585342 473854
rect 585578 473618 585662 473854
rect 585898 473618 585930 473854
rect 585310 473534 585930 473618
rect 585310 473298 585342 473534
rect 585578 473298 585662 473534
rect 585898 473298 585930 473534
rect 585310 437854 585930 473298
rect 585310 437618 585342 437854
rect 585578 437618 585662 437854
rect 585898 437618 585930 437854
rect 585310 437534 585930 437618
rect 585310 437298 585342 437534
rect 585578 437298 585662 437534
rect 585898 437298 585930 437534
rect 585310 401854 585930 437298
rect 585310 401618 585342 401854
rect 585578 401618 585662 401854
rect 585898 401618 585930 401854
rect 585310 401534 585930 401618
rect 585310 401298 585342 401534
rect 585578 401298 585662 401534
rect 585898 401298 585930 401534
rect 585310 365854 585930 401298
rect 585310 365618 585342 365854
rect 585578 365618 585662 365854
rect 585898 365618 585930 365854
rect 585310 365534 585930 365618
rect 585310 365298 585342 365534
rect 585578 365298 585662 365534
rect 585898 365298 585930 365534
rect 585310 329854 585930 365298
rect 585310 329618 585342 329854
rect 585578 329618 585662 329854
rect 585898 329618 585930 329854
rect 585310 329534 585930 329618
rect 585310 329298 585342 329534
rect 585578 329298 585662 329534
rect 585898 329298 585930 329534
rect 585310 293854 585930 329298
rect 585310 293618 585342 293854
rect 585578 293618 585662 293854
rect 585898 293618 585930 293854
rect 585310 293534 585930 293618
rect 585310 293298 585342 293534
rect 585578 293298 585662 293534
rect 585898 293298 585930 293534
rect 585310 257854 585930 293298
rect 585310 257618 585342 257854
rect 585578 257618 585662 257854
rect 585898 257618 585930 257854
rect 585310 257534 585930 257618
rect 585310 257298 585342 257534
rect 585578 257298 585662 257534
rect 585898 257298 585930 257534
rect 585310 221854 585930 257298
rect 585310 221618 585342 221854
rect 585578 221618 585662 221854
rect 585898 221618 585930 221854
rect 585310 221534 585930 221618
rect 585310 221298 585342 221534
rect 585578 221298 585662 221534
rect 585898 221298 585930 221534
rect 585310 185854 585930 221298
rect 585310 185618 585342 185854
rect 585578 185618 585662 185854
rect 585898 185618 585930 185854
rect 585310 185534 585930 185618
rect 585310 185298 585342 185534
rect 585578 185298 585662 185534
rect 585898 185298 585930 185534
rect 585310 149854 585930 185298
rect 585310 149618 585342 149854
rect 585578 149618 585662 149854
rect 585898 149618 585930 149854
rect 585310 149534 585930 149618
rect 585310 149298 585342 149534
rect 585578 149298 585662 149534
rect 585898 149298 585930 149534
rect 585310 113854 585930 149298
rect 585310 113618 585342 113854
rect 585578 113618 585662 113854
rect 585898 113618 585930 113854
rect 585310 113534 585930 113618
rect 585310 113298 585342 113534
rect 585578 113298 585662 113534
rect 585898 113298 585930 113534
rect 585310 77854 585930 113298
rect 585310 77618 585342 77854
rect 585578 77618 585662 77854
rect 585898 77618 585930 77854
rect 585310 77534 585930 77618
rect 585310 77298 585342 77534
rect 585578 77298 585662 77534
rect 585898 77298 585930 77534
rect 585310 41854 585930 77298
rect 585310 41618 585342 41854
rect 585578 41618 585662 41854
rect 585898 41618 585930 41854
rect 585310 41534 585930 41618
rect 585310 41298 585342 41534
rect 585578 41298 585662 41534
rect 585898 41298 585930 41534
rect 585310 5854 585930 41298
rect 585310 5618 585342 5854
rect 585578 5618 585662 5854
rect 585898 5618 585930 5854
rect 585310 5534 585930 5618
rect 585310 5298 585342 5534
rect 585578 5298 585662 5534
rect 585898 5298 585930 5534
rect 585310 -346 585930 5298
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 694354 586890 705242
rect 586270 694118 586302 694354
rect 586538 694118 586622 694354
rect 586858 694118 586890 694354
rect 586270 694034 586890 694118
rect 586270 693798 586302 694034
rect 586538 693798 586622 694034
rect 586858 693798 586890 694034
rect 586270 658354 586890 693798
rect 586270 658118 586302 658354
rect 586538 658118 586622 658354
rect 586858 658118 586890 658354
rect 586270 658034 586890 658118
rect 586270 657798 586302 658034
rect 586538 657798 586622 658034
rect 586858 657798 586890 658034
rect 586270 622354 586890 657798
rect 586270 622118 586302 622354
rect 586538 622118 586622 622354
rect 586858 622118 586890 622354
rect 586270 622034 586890 622118
rect 586270 621798 586302 622034
rect 586538 621798 586622 622034
rect 586858 621798 586890 622034
rect 586270 586354 586890 621798
rect 586270 586118 586302 586354
rect 586538 586118 586622 586354
rect 586858 586118 586890 586354
rect 586270 586034 586890 586118
rect 586270 585798 586302 586034
rect 586538 585798 586622 586034
rect 586858 585798 586890 586034
rect 586270 550354 586890 585798
rect 586270 550118 586302 550354
rect 586538 550118 586622 550354
rect 586858 550118 586890 550354
rect 586270 550034 586890 550118
rect 586270 549798 586302 550034
rect 586538 549798 586622 550034
rect 586858 549798 586890 550034
rect 586270 514354 586890 549798
rect 586270 514118 586302 514354
rect 586538 514118 586622 514354
rect 586858 514118 586890 514354
rect 586270 514034 586890 514118
rect 586270 513798 586302 514034
rect 586538 513798 586622 514034
rect 586858 513798 586890 514034
rect 586270 478354 586890 513798
rect 586270 478118 586302 478354
rect 586538 478118 586622 478354
rect 586858 478118 586890 478354
rect 586270 478034 586890 478118
rect 586270 477798 586302 478034
rect 586538 477798 586622 478034
rect 586858 477798 586890 478034
rect 586270 442354 586890 477798
rect 586270 442118 586302 442354
rect 586538 442118 586622 442354
rect 586858 442118 586890 442354
rect 586270 442034 586890 442118
rect 586270 441798 586302 442034
rect 586538 441798 586622 442034
rect 586858 441798 586890 442034
rect 586270 406354 586890 441798
rect 586270 406118 586302 406354
rect 586538 406118 586622 406354
rect 586858 406118 586890 406354
rect 586270 406034 586890 406118
rect 586270 405798 586302 406034
rect 586538 405798 586622 406034
rect 586858 405798 586890 406034
rect 586270 370354 586890 405798
rect 586270 370118 586302 370354
rect 586538 370118 586622 370354
rect 586858 370118 586890 370354
rect 586270 370034 586890 370118
rect 586270 369798 586302 370034
rect 586538 369798 586622 370034
rect 586858 369798 586890 370034
rect 586270 334354 586890 369798
rect 586270 334118 586302 334354
rect 586538 334118 586622 334354
rect 586858 334118 586890 334354
rect 586270 334034 586890 334118
rect 586270 333798 586302 334034
rect 586538 333798 586622 334034
rect 586858 333798 586890 334034
rect 586270 298354 586890 333798
rect 586270 298118 586302 298354
rect 586538 298118 586622 298354
rect 586858 298118 586890 298354
rect 586270 298034 586890 298118
rect 586270 297798 586302 298034
rect 586538 297798 586622 298034
rect 586858 297798 586890 298034
rect 586270 262354 586890 297798
rect 586270 262118 586302 262354
rect 586538 262118 586622 262354
rect 586858 262118 586890 262354
rect 586270 262034 586890 262118
rect 586270 261798 586302 262034
rect 586538 261798 586622 262034
rect 586858 261798 586890 262034
rect 586270 226354 586890 261798
rect 586270 226118 586302 226354
rect 586538 226118 586622 226354
rect 586858 226118 586890 226354
rect 586270 226034 586890 226118
rect 586270 225798 586302 226034
rect 586538 225798 586622 226034
rect 586858 225798 586890 226034
rect 586270 190354 586890 225798
rect 586270 190118 586302 190354
rect 586538 190118 586622 190354
rect 586858 190118 586890 190354
rect 586270 190034 586890 190118
rect 586270 189798 586302 190034
rect 586538 189798 586622 190034
rect 586858 189798 586890 190034
rect 586270 154354 586890 189798
rect 586270 154118 586302 154354
rect 586538 154118 586622 154354
rect 586858 154118 586890 154354
rect 586270 154034 586890 154118
rect 586270 153798 586302 154034
rect 586538 153798 586622 154034
rect 586858 153798 586890 154034
rect 586270 118354 586890 153798
rect 586270 118118 586302 118354
rect 586538 118118 586622 118354
rect 586858 118118 586890 118354
rect 586270 118034 586890 118118
rect 586270 117798 586302 118034
rect 586538 117798 586622 118034
rect 586858 117798 586890 118034
rect 586270 82354 586890 117798
rect 586270 82118 586302 82354
rect 586538 82118 586622 82354
rect 586858 82118 586890 82354
rect 586270 82034 586890 82118
rect 586270 81798 586302 82034
rect 586538 81798 586622 82034
rect 586858 81798 586890 82034
rect 586270 46354 586890 81798
rect 586270 46118 586302 46354
rect 586538 46118 586622 46354
rect 586858 46118 586890 46354
rect 586270 46034 586890 46118
rect 586270 45798 586302 46034
rect 586538 45798 586622 46034
rect 586858 45798 586890 46034
rect 586270 10354 586890 45798
rect 586270 10118 586302 10354
rect 586538 10118 586622 10354
rect 586858 10118 586890 10354
rect 586270 10034 586890 10118
rect 586270 9798 586302 10034
rect 586538 9798 586622 10034
rect 586858 9798 586890 10034
rect 582294 -1542 582326 -1306
rect 582562 -1542 582646 -1306
rect 582882 -1542 582914 -1306
rect 582294 -1626 582914 -1542
rect 582294 -1862 582326 -1626
rect 582562 -1862 582646 -1626
rect 582882 -1862 582914 -1626
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 582294 -7654 582914 -1862
rect 586270 -1306 586890 9798
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 -2266 587850 706202
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 -3226 588810 707162
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 -4186 589770 708122
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 -5146 590730 709082
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 -6106 591690 710042
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 -7066 592650 711002
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 582326 705562 582562 705798
rect 582646 705562 582882 705798
rect 582326 705242 582562 705478
rect 582646 705242 582882 705478
rect -2934 694118 -2698 694354
rect -2614 694118 -2378 694354
rect -2934 693798 -2698 694034
rect -2614 693798 -2378 694034
rect -2934 658118 -2698 658354
rect -2614 658118 -2378 658354
rect -2934 657798 -2698 658034
rect -2614 657798 -2378 658034
rect -2934 622118 -2698 622354
rect -2614 622118 -2378 622354
rect -2934 621798 -2698 622034
rect -2614 621798 -2378 622034
rect -2934 586118 -2698 586354
rect -2614 586118 -2378 586354
rect -2934 585798 -2698 586034
rect -2614 585798 -2378 586034
rect -2934 550118 -2698 550354
rect -2614 550118 -2378 550354
rect -2934 549798 -2698 550034
rect -2614 549798 -2378 550034
rect -2934 514118 -2698 514354
rect -2614 514118 -2378 514354
rect -2934 513798 -2698 514034
rect -2614 513798 -2378 514034
rect -2934 478118 -2698 478354
rect -2614 478118 -2378 478354
rect -2934 477798 -2698 478034
rect -2614 477798 -2378 478034
rect -2934 442118 -2698 442354
rect -2614 442118 -2378 442354
rect -2934 441798 -2698 442034
rect -2614 441798 -2378 442034
rect -2934 406118 -2698 406354
rect -2614 406118 -2378 406354
rect -2934 405798 -2698 406034
rect -2614 405798 -2378 406034
rect -2934 370118 -2698 370354
rect -2614 370118 -2378 370354
rect -2934 369798 -2698 370034
rect -2614 369798 -2378 370034
rect -2934 334118 -2698 334354
rect -2614 334118 -2378 334354
rect -2934 333798 -2698 334034
rect -2614 333798 -2378 334034
rect -2934 298118 -2698 298354
rect -2614 298118 -2378 298354
rect -2934 297798 -2698 298034
rect -2614 297798 -2378 298034
rect -2934 262118 -2698 262354
rect -2614 262118 -2378 262354
rect -2934 261798 -2698 262034
rect -2614 261798 -2378 262034
rect -2934 226118 -2698 226354
rect -2614 226118 -2378 226354
rect -2934 225798 -2698 226034
rect -2614 225798 -2378 226034
rect -2934 190118 -2698 190354
rect -2614 190118 -2378 190354
rect -2934 189798 -2698 190034
rect -2614 189798 -2378 190034
rect -2934 154118 -2698 154354
rect -2614 154118 -2378 154354
rect -2934 153798 -2698 154034
rect -2614 153798 -2378 154034
rect -2934 118118 -2698 118354
rect -2614 118118 -2378 118354
rect -2934 117798 -2698 118034
rect -2614 117798 -2378 118034
rect -2934 82118 -2698 82354
rect -2614 82118 -2378 82354
rect -2934 81798 -2698 82034
rect -2614 81798 -2378 82034
rect -2934 46118 -2698 46354
rect -2614 46118 -2378 46354
rect -2934 45798 -2698 46034
rect -2614 45798 -2378 46034
rect -2934 10118 -2698 10354
rect -2614 10118 -2378 10354
rect -2934 9798 -2698 10034
rect -2614 9798 -2378 10034
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 23826 694118 24062 694354
rect 24146 694118 24382 694354
rect 23826 693798 24062 694034
rect 24146 693798 24382 694034
rect 59826 694118 60062 694354
rect 60146 694118 60382 694354
rect 59826 693798 60062 694034
rect 60146 693798 60382 694034
rect 95826 694118 96062 694354
rect 96146 694118 96382 694354
rect 95826 693798 96062 694034
rect 96146 693798 96382 694034
rect 131826 694118 132062 694354
rect 132146 694118 132382 694354
rect 131826 693798 132062 694034
rect 132146 693798 132382 694034
rect 167826 694118 168062 694354
rect 168146 694118 168382 694354
rect 167826 693798 168062 694034
rect 168146 693798 168382 694034
rect 203826 694118 204062 694354
rect 204146 694118 204382 694354
rect 203826 693798 204062 694034
rect 204146 693798 204382 694034
rect 239826 694118 240062 694354
rect 240146 694118 240382 694354
rect 239826 693798 240062 694034
rect 240146 693798 240382 694034
rect 275826 694118 276062 694354
rect 276146 694118 276382 694354
rect 275826 693798 276062 694034
rect 276146 693798 276382 694034
rect 311826 694118 312062 694354
rect 312146 694118 312382 694354
rect 311826 693798 312062 694034
rect 312146 693798 312382 694034
rect 347826 694118 348062 694354
rect 348146 694118 348382 694354
rect 347826 693798 348062 694034
rect 348146 693798 348382 694034
rect 383826 694118 384062 694354
rect 384146 694118 384382 694354
rect 383826 693798 384062 694034
rect 384146 693798 384382 694034
rect 419826 694118 420062 694354
rect 420146 694118 420382 694354
rect 419826 693798 420062 694034
rect 420146 693798 420382 694034
rect 455826 694118 456062 694354
rect 456146 694118 456382 694354
rect 455826 693798 456062 694034
rect 456146 693798 456382 694034
rect 491826 694118 492062 694354
rect 492146 694118 492382 694354
rect 491826 693798 492062 694034
rect 492146 693798 492382 694034
rect 527826 694118 528062 694354
rect 528146 694118 528382 694354
rect 527826 693798 528062 694034
rect 528146 693798 528382 694034
rect 563826 694118 564062 694354
rect 564146 694118 564382 694354
rect 563826 693798 564062 694034
rect 564146 693798 564382 694034
rect 582326 694118 582562 694354
rect 582646 694118 582882 694354
rect 582326 693798 582562 694034
rect 582646 693798 582882 694034
rect -1974 689618 -1738 689854
rect -1654 689618 -1418 689854
rect -1974 689298 -1738 689534
rect -1654 689298 -1418 689534
rect 5826 689618 6062 689854
rect 6146 689618 6382 689854
rect 5826 689298 6062 689534
rect 6146 689298 6382 689534
rect 41826 689618 42062 689854
rect 42146 689618 42382 689854
rect 41826 689298 42062 689534
rect 42146 689298 42382 689534
rect 77826 689618 78062 689854
rect 78146 689618 78382 689854
rect 77826 689298 78062 689534
rect 78146 689298 78382 689534
rect 113826 689618 114062 689854
rect 114146 689618 114382 689854
rect 113826 689298 114062 689534
rect 114146 689298 114382 689534
rect 149826 689618 150062 689854
rect 150146 689618 150382 689854
rect 149826 689298 150062 689534
rect 150146 689298 150382 689534
rect 185826 689618 186062 689854
rect 186146 689618 186382 689854
rect 185826 689298 186062 689534
rect 186146 689298 186382 689534
rect 221826 689618 222062 689854
rect 222146 689618 222382 689854
rect 221826 689298 222062 689534
rect 222146 689298 222382 689534
rect 257826 689618 258062 689854
rect 258146 689618 258382 689854
rect 257826 689298 258062 689534
rect 258146 689298 258382 689534
rect 293826 689618 294062 689854
rect 294146 689618 294382 689854
rect 293826 689298 294062 689534
rect 294146 689298 294382 689534
rect 329826 689618 330062 689854
rect 330146 689618 330382 689854
rect 329826 689298 330062 689534
rect 330146 689298 330382 689534
rect 365826 689618 366062 689854
rect 366146 689618 366382 689854
rect 365826 689298 366062 689534
rect 366146 689298 366382 689534
rect 401826 689618 402062 689854
rect 402146 689618 402382 689854
rect 401826 689298 402062 689534
rect 402146 689298 402382 689534
rect 437826 689618 438062 689854
rect 438146 689618 438382 689854
rect 437826 689298 438062 689534
rect 438146 689298 438382 689534
rect 473826 689618 474062 689854
rect 474146 689618 474382 689854
rect 473826 689298 474062 689534
rect 474146 689298 474382 689534
rect 509826 689618 510062 689854
rect 510146 689618 510382 689854
rect 509826 689298 510062 689534
rect 510146 689298 510382 689534
rect 545826 689618 546062 689854
rect 546146 689618 546382 689854
rect 545826 689298 546062 689534
rect 546146 689298 546382 689534
rect 13198 658118 13434 658354
rect 13518 658118 13754 658354
rect 13198 657798 13434 658034
rect 13518 657798 13754 658034
rect 167826 658118 168062 658354
rect 168146 658118 168382 658354
rect 167826 657798 168062 658034
rect 168146 657798 168382 658034
rect 291590 658118 291826 658354
rect 291910 658118 292146 658354
rect 291590 657798 291826 658034
rect 291910 657798 292146 658034
rect 419826 658118 420062 658354
rect 420146 658118 420382 658354
rect 419826 657798 420062 658034
rect 420146 657798 420382 658034
rect 563826 658118 564062 658354
rect 564146 658118 564382 658354
rect 563826 657798 564062 658034
rect 564146 657798 564382 658034
rect 582326 658118 582562 658354
rect 582646 658118 582882 658354
rect 582326 657798 582562 658034
rect 582646 657798 582882 658034
rect -1974 653618 -1738 653854
rect -1654 653618 -1418 653854
rect -1974 653298 -1738 653534
rect -1654 653298 -1418 653534
rect 5826 653618 6062 653854
rect 6146 653618 6382 653854
rect 5826 653298 6062 653534
rect 6146 653298 6382 653534
rect 173094 653618 173330 653854
rect 173414 653618 173650 653854
rect 173094 653298 173330 653534
rect 173414 653298 173650 653534
rect 293826 653618 294062 653854
rect 294146 653618 294382 653854
rect 293826 653298 294062 653534
rect 294146 653298 294382 653534
rect 401826 653618 402062 653854
rect 402146 653618 402382 653854
rect 401826 653298 402062 653534
rect 402146 653298 402382 653534
rect 570350 653618 570586 653854
rect 570670 653618 570906 653854
rect 570350 653298 570586 653534
rect 570670 653298 570906 653534
rect 13198 622118 13434 622354
rect 13518 622118 13754 622354
rect 13198 621798 13434 622034
rect 13518 621798 13754 622034
rect 167826 622118 168062 622354
rect 168146 622118 168382 622354
rect 167826 621798 168062 622034
rect 168146 621798 168382 622034
rect 291590 622118 291826 622354
rect 291910 622118 292146 622354
rect 291590 621798 291826 622034
rect 291910 621798 292146 622034
rect 419826 622118 420062 622354
rect 420146 622118 420382 622354
rect 419826 621798 420062 622034
rect 420146 621798 420382 622034
rect 563826 622118 564062 622354
rect 564146 622118 564382 622354
rect 563826 621798 564062 622034
rect 564146 621798 564382 622034
rect 582326 622118 582562 622354
rect 582646 622118 582882 622354
rect 582326 621798 582562 622034
rect 582646 621798 582882 622034
rect -1974 617618 -1738 617854
rect -1654 617618 -1418 617854
rect -1974 617298 -1738 617534
rect -1654 617298 -1418 617534
rect 5826 617618 6062 617854
rect 6146 617618 6382 617854
rect 5826 617298 6062 617534
rect 6146 617298 6382 617534
rect 173094 617618 173330 617854
rect 173414 617618 173650 617854
rect 173094 617298 173330 617534
rect 173414 617298 173650 617534
rect 293826 617618 294062 617854
rect 294146 617618 294382 617854
rect 293826 617298 294062 617534
rect 294146 617298 294382 617534
rect 401826 617618 402062 617854
rect 402146 617618 402382 617854
rect 401826 617298 402062 617534
rect 402146 617298 402382 617534
rect 570350 617618 570586 617854
rect 570670 617618 570906 617854
rect 570350 617298 570586 617534
rect 570670 617298 570906 617534
rect 23826 586118 24062 586354
rect 24146 586118 24382 586354
rect 23826 585798 24062 586034
rect 24146 585798 24382 586034
rect 59826 586118 60062 586354
rect 60146 586118 60382 586354
rect 59826 585798 60062 586034
rect 60146 585798 60382 586034
rect 95826 586118 96062 586354
rect 96146 586118 96382 586354
rect 95826 585798 96062 586034
rect 96146 585798 96382 586034
rect 131826 586118 132062 586354
rect 132146 586118 132382 586354
rect 131826 585798 132062 586034
rect 132146 585798 132382 586034
rect 167826 586118 168062 586354
rect 168146 586118 168382 586354
rect 167826 585798 168062 586034
rect 168146 585798 168382 586034
rect 203826 586118 204062 586354
rect 204146 586118 204382 586354
rect 203826 585798 204062 586034
rect 204146 585798 204382 586034
rect 239826 586118 240062 586354
rect 240146 586118 240382 586354
rect 239826 585798 240062 586034
rect 240146 585798 240382 586034
rect 275826 586118 276062 586354
rect 276146 586118 276382 586354
rect 275826 585798 276062 586034
rect 276146 585798 276382 586034
rect 311826 586118 312062 586354
rect 312146 586118 312382 586354
rect 311826 585798 312062 586034
rect 312146 585798 312382 586034
rect 347826 586118 348062 586354
rect 348146 586118 348382 586354
rect 347826 585798 348062 586034
rect 348146 585798 348382 586034
rect 383826 586118 384062 586354
rect 384146 586118 384382 586354
rect 383826 585798 384062 586034
rect 384146 585798 384382 586034
rect 419826 586118 420062 586354
rect 420146 586118 420382 586354
rect 419826 585798 420062 586034
rect 420146 585798 420382 586034
rect 455826 586118 456062 586354
rect 456146 586118 456382 586354
rect 455826 585798 456062 586034
rect 456146 585798 456382 586034
rect 491826 586118 492062 586354
rect 492146 586118 492382 586354
rect 491826 585798 492062 586034
rect 492146 585798 492382 586034
rect 527826 586118 528062 586354
rect 528146 586118 528382 586354
rect 527826 585798 528062 586034
rect 528146 585798 528382 586034
rect 563826 586118 564062 586354
rect 564146 586118 564382 586354
rect 563826 585798 564062 586034
rect 564146 585798 564382 586034
rect 582326 586118 582562 586354
rect 582646 586118 582882 586354
rect 582326 585798 582562 586034
rect 582646 585798 582882 586034
rect -1974 581618 -1738 581854
rect -1654 581618 -1418 581854
rect -1974 581298 -1738 581534
rect -1654 581298 -1418 581534
rect 5826 581618 6062 581854
rect 6146 581618 6382 581854
rect 5826 581298 6062 581534
rect 6146 581298 6382 581534
rect 41826 581618 42062 581854
rect 42146 581618 42382 581854
rect 41826 581298 42062 581534
rect 42146 581298 42382 581534
rect 77826 581618 78062 581854
rect 78146 581618 78382 581854
rect 77826 581298 78062 581534
rect 78146 581298 78382 581534
rect 113826 581618 114062 581854
rect 114146 581618 114382 581854
rect 113826 581298 114062 581534
rect 114146 581298 114382 581534
rect 149826 581618 150062 581854
rect 150146 581618 150382 581854
rect 149826 581298 150062 581534
rect 150146 581298 150382 581534
rect 185826 581618 186062 581854
rect 186146 581618 186382 581854
rect 185826 581298 186062 581534
rect 186146 581298 186382 581534
rect 221826 581618 222062 581854
rect 222146 581618 222382 581854
rect 221826 581298 222062 581534
rect 222146 581298 222382 581534
rect 257826 581618 258062 581854
rect 258146 581618 258382 581854
rect 257826 581298 258062 581534
rect 258146 581298 258382 581534
rect 293826 581618 294062 581854
rect 294146 581618 294382 581854
rect 293826 581298 294062 581534
rect 294146 581298 294382 581534
rect 329826 581618 330062 581854
rect 330146 581618 330382 581854
rect 329826 581298 330062 581534
rect 330146 581298 330382 581534
rect 365826 581618 366062 581854
rect 366146 581618 366382 581854
rect 365826 581298 366062 581534
rect 366146 581298 366382 581534
rect 401826 581618 402062 581854
rect 402146 581618 402382 581854
rect 401826 581298 402062 581534
rect 402146 581298 402382 581534
rect 437826 581618 438062 581854
rect 438146 581618 438382 581854
rect 437826 581298 438062 581534
rect 438146 581298 438382 581534
rect 473826 581618 474062 581854
rect 474146 581618 474382 581854
rect 473826 581298 474062 581534
rect 474146 581298 474382 581534
rect 509826 581618 510062 581854
rect 510146 581618 510382 581854
rect 509826 581298 510062 581534
rect 510146 581298 510382 581534
rect 545826 581618 546062 581854
rect 546146 581618 546382 581854
rect 545826 581298 546062 581534
rect 546146 581298 546382 581534
rect 13198 550118 13434 550354
rect 13518 550118 13754 550354
rect 13198 549798 13434 550034
rect 13518 549798 13754 550034
rect 167826 550118 168062 550354
rect 168146 550118 168382 550354
rect 167826 549798 168062 550034
rect 168146 549798 168382 550034
rect 203826 550118 204062 550354
rect 204146 550118 204382 550354
rect 203826 549798 204062 550034
rect 204146 549798 204382 550034
rect 239826 550118 240062 550354
rect 240146 550118 240382 550354
rect 239826 549798 240062 550034
rect 240146 549798 240382 550034
rect 275826 550118 276062 550354
rect 276146 550118 276382 550354
rect 275826 549798 276062 550034
rect 276146 549798 276382 550034
rect 311826 550118 312062 550354
rect 312146 550118 312382 550354
rect 311826 549798 312062 550034
rect 312146 549798 312382 550034
rect 347826 550118 348062 550354
rect 348146 550118 348382 550354
rect 347826 549798 348062 550034
rect 348146 549798 348382 550034
rect 383826 550118 384062 550354
rect 384146 550118 384382 550354
rect 383826 549798 384062 550034
rect 384146 549798 384382 550034
rect 419826 550118 420062 550354
rect 420146 550118 420382 550354
rect 419826 549798 420062 550034
rect 420146 549798 420382 550034
rect 563826 550118 564062 550354
rect 564146 550118 564382 550354
rect 563826 549798 564062 550034
rect 564146 549798 564382 550034
rect 582326 550118 582562 550354
rect 582646 550118 582882 550354
rect 582326 549798 582562 550034
rect 582646 549798 582882 550034
rect -1974 545618 -1738 545854
rect -1654 545618 -1418 545854
rect -1974 545298 -1738 545534
rect -1654 545298 -1418 545534
rect 5826 545618 6062 545854
rect 6146 545618 6382 545854
rect 5826 545298 6062 545534
rect 6146 545298 6382 545534
rect 185826 545618 186062 545854
rect 186146 545618 186382 545854
rect 185826 545298 186062 545534
rect 186146 545298 186382 545534
rect 221826 545618 222062 545854
rect 222146 545618 222382 545854
rect 221826 545298 222062 545534
rect 222146 545298 222382 545534
rect 257826 545618 258062 545854
rect 258146 545618 258382 545854
rect 257826 545298 258062 545534
rect 258146 545298 258382 545534
rect 293826 545618 294062 545854
rect 294146 545618 294382 545854
rect 293826 545298 294062 545534
rect 294146 545298 294382 545534
rect 329826 545618 330062 545854
rect 330146 545618 330382 545854
rect 329826 545298 330062 545534
rect 330146 545298 330382 545534
rect 365826 545618 366062 545854
rect 366146 545618 366382 545854
rect 365826 545298 366062 545534
rect 366146 545298 366382 545534
rect 401826 545618 402062 545854
rect 402146 545618 402382 545854
rect 401826 545298 402062 545534
rect 402146 545298 402382 545534
rect 570350 545618 570586 545854
rect 570670 545618 570906 545854
rect 570350 545298 570586 545534
rect 570670 545298 570906 545534
rect 13198 514118 13434 514354
rect 13518 514118 13754 514354
rect 13198 513798 13434 514034
rect 13518 513798 13754 514034
rect 167826 514118 168062 514354
rect 168146 514118 168382 514354
rect 167826 513798 168062 514034
rect 168146 513798 168382 514034
rect 203826 514118 204062 514354
rect 204146 514118 204382 514354
rect 203826 513798 204062 514034
rect 204146 513798 204382 514034
rect 239826 514118 240062 514354
rect 240146 514118 240382 514354
rect 239826 513798 240062 514034
rect 240146 513798 240382 514034
rect 275826 514118 276062 514354
rect 276146 514118 276382 514354
rect 275826 513798 276062 514034
rect 276146 513798 276382 514034
rect 311826 514118 312062 514354
rect 312146 514118 312382 514354
rect 311826 513798 312062 514034
rect 312146 513798 312382 514034
rect 347826 514118 348062 514354
rect 348146 514118 348382 514354
rect 347826 513798 348062 514034
rect 348146 513798 348382 514034
rect 383826 514118 384062 514354
rect 384146 514118 384382 514354
rect 383826 513798 384062 514034
rect 384146 513798 384382 514034
rect 419826 514118 420062 514354
rect 420146 514118 420382 514354
rect 419826 513798 420062 514034
rect 420146 513798 420382 514034
rect 563826 514118 564062 514354
rect 564146 514118 564382 514354
rect 563826 513798 564062 514034
rect 564146 513798 564382 514034
rect 582326 514118 582562 514354
rect 582646 514118 582882 514354
rect 582326 513798 582562 514034
rect 582646 513798 582882 514034
rect -1974 509618 -1738 509854
rect -1654 509618 -1418 509854
rect -1974 509298 -1738 509534
rect -1654 509298 -1418 509534
rect 5826 509618 6062 509854
rect 6146 509618 6382 509854
rect 5826 509298 6062 509534
rect 6146 509298 6382 509534
rect 185826 509618 186062 509854
rect 186146 509618 186382 509854
rect 185826 509298 186062 509534
rect 186146 509298 186382 509534
rect 221826 509618 222062 509854
rect 222146 509618 222382 509854
rect 221826 509298 222062 509534
rect 222146 509298 222382 509534
rect 257826 509618 258062 509854
rect 258146 509618 258382 509854
rect 257826 509298 258062 509534
rect 258146 509298 258382 509534
rect 293826 509618 294062 509854
rect 294146 509618 294382 509854
rect 293826 509298 294062 509534
rect 294146 509298 294382 509534
rect 329826 509618 330062 509854
rect 330146 509618 330382 509854
rect 329826 509298 330062 509534
rect 330146 509298 330382 509534
rect 365826 509618 366062 509854
rect 366146 509618 366382 509854
rect 365826 509298 366062 509534
rect 366146 509298 366382 509534
rect 401826 509618 402062 509854
rect 402146 509618 402382 509854
rect 401826 509298 402062 509534
rect 402146 509298 402382 509534
rect 570350 509618 570586 509854
rect 570670 509618 570906 509854
rect 570350 509298 570586 509534
rect 570670 509298 570906 509534
rect 23826 478118 24062 478354
rect 24146 478118 24382 478354
rect 23826 477798 24062 478034
rect 24146 477798 24382 478034
rect 59826 478118 60062 478354
rect 60146 478118 60382 478354
rect 59826 477798 60062 478034
rect 60146 477798 60382 478034
rect 95826 478118 96062 478354
rect 96146 478118 96382 478354
rect 95826 477798 96062 478034
rect 96146 477798 96382 478034
rect 131826 478118 132062 478354
rect 132146 478118 132382 478354
rect 131826 477798 132062 478034
rect 132146 477798 132382 478034
rect 167826 478118 168062 478354
rect 168146 478118 168382 478354
rect 167826 477798 168062 478034
rect 168146 477798 168382 478034
rect 203826 478118 204062 478354
rect 204146 478118 204382 478354
rect 203826 477798 204062 478034
rect 204146 477798 204382 478034
rect 239826 478118 240062 478354
rect 240146 478118 240382 478354
rect 239826 477798 240062 478034
rect 240146 477798 240382 478034
rect 275826 478118 276062 478354
rect 276146 478118 276382 478354
rect 275826 477798 276062 478034
rect 276146 477798 276382 478034
rect 311826 478118 312062 478354
rect 312146 478118 312382 478354
rect 311826 477798 312062 478034
rect 312146 477798 312382 478034
rect 347826 478118 348062 478354
rect 348146 478118 348382 478354
rect 347826 477798 348062 478034
rect 348146 477798 348382 478034
rect 383826 478118 384062 478354
rect 384146 478118 384382 478354
rect 383826 477798 384062 478034
rect 384146 477798 384382 478034
rect 419826 478118 420062 478354
rect 420146 478118 420382 478354
rect 419826 477798 420062 478034
rect 420146 477798 420382 478034
rect 455826 478118 456062 478354
rect 456146 478118 456382 478354
rect 455826 477798 456062 478034
rect 456146 477798 456382 478034
rect 491826 478118 492062 478354
rect 492146 478118 492382 478354
rect 491826 477798 492062 478034
rect 492146 477798 492382 478034
rect 527826 478118 528062 478354
rect 528146 478118 528382 478354
rect 527826 477798 528062 478034
rect 528146 477798 528382 478034
rect 563826 478118 564062 478354
rect 564146 478118 564382 478354
rect 563826 477798 564062 478034
rect 564146 477798 564382 478034
rect 582326 478118 582562 478354
rect 582646 478118 582882 478354
rect 582326 477798 582562 478034
rect 582646 477798 582882 478034
rect -1974 473618 -1738 473854
rect -1654 473618 -1418 473854
rect -1974 473298 -1738 473534
rect -1654 473298 -1418 473534
rect 5826 473618 6062 473854
rect 6146 473618 6382 473854
rect 5826 473298 6062 473534
rect 6146 473298 6382 473534
rect 41826 473618 42062 473854
rect 42146 473618 42382 473854
rect 41826 473298 42062 473534
rect 42146 473298 42382 473534
rect 77826 473618 78062 473854
rect 78146 473618 78382 473854
rect 77826 473298 78062 473534
rect 78146 473298 78382 473534
rect 113826 473618 114062 473854
rect 114146 473618 114382 473854
rect 113826 473298 114062 473534
rect 114146 473298 114382 473534
rect 149826 473618 150062 473854
rect 150146 473618 150382 473854
rect 149826 473298 150062 473534
rect 150146 473298 150382 473534
rect 185826 473618 186062 473854
rect 186146 473618 186382 473854
rect 185826 473298 186062 473534
rect 186146 473298 186382 473534
rect 221826 473618 222062 473854
rect 222146 473618 222382 473854
rect 221826 473298 222062 473534
rect 222146 473298 222382 473534
rect 257826 473618 258062 473854
rect 258146 473618 258382 473854
rect 257826 473298 258062 473534
rect 258146 473298 258382 473534
rect 293826 473618 294062 473854
rect 294146 473618 294382 473854
rect 293826 473298 294062 473534
rect 294146 473298 294382 473534
rect 329826 473618 330062 473854
rect 330146 473618 330382 473854
rect 329826 473298 330062 473534
rect 330146 473298 330382 473534
rect 365826 473618 366062 473854
rect 366146 473618 366382 473854
rect 365826 473298 366062 473534
rect 366146 473298 366382 473534
rect 401826 473618 402062 473854
rect 402146 473618 402382 473854
rect 401826 473298 402062 473534
rect 402146 473298 402382 473534
rect 437826 473618 438062 473854
rect 438146 473618 438382 473854
rect 437826 473298 438062 473534
rect 438146 473298 438382 473534
rect 473826 473618 474062 473854
rect 474146 473618 474382 473854
rect 473826 473298 474062 473534
rect 474146 473298 474382 473534
rect 509826 473618 510062 473854
rect 510146 473618 510382 473854
rect 509826 473298 510062 473534
rect 510146 473298 510382 473534
rect 545826 473618 546062 473854
rect 546146 473618 546382 473854
rect 545826 473298 546062 473534
rect 546146 473298 546382 473534
rect 13198 442118 13434 442354
rect 13518 442118 13754 442354
rect 13198 441798 13434 442034
rect 13518 441798 13754 442034
rect 167826 442118 168062 442354
rect 168146 442118 168382 442354
rect 167826 441798 168062 442034
rect 168146 441798 168382 442034
rect 203826 442118 204062 442354
rect 204146 442118 204382 442354
rect 203826 441798 204062 442034
rect 204146 441798 204382 442034
rect 239826 442118 240062 442354
rect 240146 442118 240382 442354
rect 239826 441798 240062 442034
rect 240146 441798 240382 442034
rect 275826 442118 276062 442354
rect 276146 442118 276382 442354
rect 275826 441798 276062 442034
rect 276146 441798 276382 442034
rect 311826 442118 312062 442354
rect 312146 442118 312382 442354
rect 311826 441798 312062 442034
rect 312146 441798 312382 442034
rect 347826 442118 348062 442354
rect 348146 442118 348382 442354
rect 347826 441798 348062 442034
rect 348146 441798 348382 442034
rect 383826 442118 384062 442354
rect 384146 442118 384382 442354
rect 383826 441798 384062 442034
rect 384146 441798 384382 442034
rect 419826 442118 420062 442354
rect 420146 442118 420382 442354
rect 419826 441798 420062 442034
rect 420146 441798 420382 442034
rect 563826 442118 564062 442354
rect 564146 442118 564382 442354
rect 563826 441798 564062 442034
rect 564146 441798 564382 442034
rect 582326 442118 582562 442354
rect 582646 442118 582882 442354
rect 582326 441798 582562 442034
rect 582646 441798 582882 442034
rect -1974 437618 -1738 437854
rect -1654 437618 -1418 437854
rect -1974 437298 -1738 437534
rect -1654 437298 -1418 437534
rect 5826 437618 6062 437854
rect 6146 437618 6382 437854
rect 5826 437298 6062 437534
rect 6146 437298 6382 437534
rect 185826 437618 186062 437854
rect 186146 437618 186382 437854
rect 185826 437298 186062 437534
rect 186146 437298 186382 437534
rect 221826 437618 222062 437854
rect 222146 437618 222382 437854
rect 221826 437298 222062 437534
rect 222146 437298 222382 437534
rect 257826 437618 258062 437854
rect 258146 437618 258382 437854
rect 257826 437298 258062 437534
rect 258146 437298 258382 437534
rect 293826 437618 294062 437854
rect 294146 437618 294382 437854
rect 293826 437298 294062 437534
rect 294146 437298 294382 437534
rect 329826 437618 330062 437854
rect 330146 437618 330382 437854
rect 329826 437298 330062 437534
rect 330146 437298 330382 437534
rect 365826 437618 366062 437854
rect 366146 437618 366382 437854
rect 365826 437298 366062 437534
rect 366146 437298 366382 437534
rect 401826 437618 402062 437854
rect 402146 437618 402382 437854
rect 401826 437298 402062 437534
rect 402146 437298 402382 437534
rect 570350 437618 570586 437854
rect 570670 437618 570906 437854
rect 570350 437298 570586 437534
rect 570670 437298 570906 437534
rect 13198 406118 13434 406354
rect 13518 406118 13754 406354
rect 13198 405798 13434 406034
rect 13518 405798 13754 406034
rect 167826 406118 168062 406354
rect 168146 406118 168382 406354
rect 167826 405798 168062 406034
rect 168146 405798 168382 406034
rect 203826 406118 204062 406354
rect 204146 406118 204382 406354
rect 203826 405798 204062 406034
rect 204146 405798 204382 406034
rect 239826 406118 240062 406354
rect 240146 406118 240382 406354
rect 239826 405798 240062 406034
rect 240146 405798 240382 406034
rect 275826 406118 276062 406354
rect 276146 406118 276382 406354
rect 275826 405798 276062 406034
rect 276146 405798 276382 406034
rect 311826 406118 312062 406354
rect 312146 406118 312382 406354
rect 311826 405798 312062 406034
rect 312146 405798 312382 406034
rect 347826 406118 348062 406354
rect 348146 406118 348382 406354
rect 347826 405798 348062 406034
rect 348146 405798 348382 406034
rect 383826 406118 384062 406354
rect 384146 406118 384382 406354
rect 383826 405798 384062 406034
rect 384146 405798 384382 406034
rect 419826 406118 420062 406354
rect 420146 406118 420382 406354
rect 419826 405798 420062 406034
rect 420146 405798 420382 406034
rect 563826 406118 564062 406354
rect 564146 406118 564382 406354
rect 563826 405798 564062 406034
rect 564146 405798 564382 406034
rect 582326 406118 582562 406354
rect 582646 406118 582882 406354
rect 582326 405798 582562 406034
rect 582646 405798 582882 406034
rect -1974 401618 -1738 401854
rect -1654 401618 -1418 401854
rect -1974 401298 -1738 401534
rect -1654 401298 -1418 401534
rect 5826 401618 6062 401854
rect 6146 401618 6382 401854
rect 5826 401298 6062 401534
rect 6146 401298 6382 401534
rect 185826 401618 186062 401854
rect 186146 401618 186382 401854
rect 185826 401298 186062 401534
rect 186146 401298 186382 401534
rect 221826 401618 222062 401854
rect 222146 401618 222382 401854
rect 221826 401298 222062 401534
rect 222146 401298 222382 401534
rect 257826 401618 258062 401854
rect 258146 401618 258382 401854
rect 257826 401298 258062 401534
rect 258146 401298 258382 401534
rect 293826 401618 294062 401854
rect 294146 401618 294382 401854
rect 293826 401298 294062 401534
rect 294146 401298 294382 401534
rect 329826 401618 330062 401854
rect 330146 401618 330382 401854
rect 329826 401298 330062 401534
rect 330146 401298 330382 401534
rect 365826 401618 366062 401854
rect 366146 401618 366382 401854
rect 365826 401298 366062 401534
rect 366146 401298 366382 401534
rect 401826 401618 402062 401854
rect 402146 401618 402382 401854
rect 401826 401298 402062 401534
rect 402146 401298 402382 401534
rect 570350 401618 570586 401854
rect 570670 401618 570906 401854
rect 570350 401298 570586 401534
rect 570670 401298 570906 401534
rect 13198 370118 13434 370354
rect 13518 370118 13754 370354
rect 13198 369798 13434 370034
rect 13518 369798 13754 370034
rect 167826 370118 168062 370354
rect 168146 370118 168382 370354
rect 167826 369798 168062 370034
rect 168146 369798 168382 370034
rect 203826 370118 204062 370354
rect 204146 370118 204382 370354
rect 203826 369798 204062 370034
rect 204146 369798 204382 370034
rect 239826 370118 240062 370354
rect 240146 370118 240382 370354
rect 239826 369798 240062 370034
rect 240146 369798 240382 370034
rect 275826 370118 276062 370354
rect 276146 370118 276382 370354
rect 275826 369798 276062 370034
rect 276146 369798 276382 370034
rect 311826 370118 312062 370354
rect 312146 370118 312382 370354
rect 311826 369798 312062 370034
rect 312146 369798 312382 370034
rect 347826 370118 348062 370354
rect 348146 370118 348382 370354
rect 347826 369798 348062 370034
rect 348146 369798 348382 370034
rect 383826 370118 384062 370354
rect 384146 370118 384382 370354
rect 383826 369798 384062 370034
rect 384146 369798 384382 370034
rect 419826 370118 420062 370354
rect 420146 370118 420382 370354
rect 419826 369798 420062 370034
rect 420146 369798 420382 370034
rect 563826 370118 564062 370354
rect 564146 370118 564382 370354
rect 563826 369798 564062 370034
rect 564146 369798 564382 370034
rect 582326 370118 582562 370354
rect 582646 370118 582882 370354
rect 582326 369798 582562 370034
rect 582646 369798 582882 370034
rect -1974 365618 -1738 365854
rect -1654 365618 -1418 365854
rect -1974 365298 -1738 365534
rect -1654 365298 -1418 365534
rect 5826 365618 6062 365854
rect 6146 365618 6382 365854
rect 5826 365298 6062 365534
rect 6146 365298 6382 365534
rect 41826 365618 42062 365854
rect 42146 365618 42382 365854
rect 41826 365298 42062 365534
rect 42146 365298 42382 365534
rect 77826 365618 78062 365854
rect 78146 365618 78382 365854
rect 77826 365298 78062 365534
rect 78146 365298 78382 365534
rect 113826 365618 114062 365854
rect 114146 365618 114382 365854
rect 113826 365298 114062 365534
rect 114146 365298 114382 365534
rect 149826 365618 150062 365854
rect 150146 365618 150382 365854
rect 149826 365298 150062 365534
rect 150146 365298 150382 365534
rect 185826 365618 186062 365854
rect 186146 365618 186382 365854
rect 185826 365298 186062 365534
rect 186146 365298 186382 365534
rect 221826 365618 222062 365854
rect 222146 365618 222382 365854
rect 221826 365298 222062 365534
rect 222146 365298 222382 365534
rect 257826 365618 258062 365854
rect 258146 365618 258382 365854
rect 257826 365298 258062 365534
rect 258146 365298 258382 365534
rect 293826 365618 294062 365854
rect 294146 365618 294382 365854
rect 293826 365298 294062 365534
rect 294146 365298 294382 365534
rect 329826 365618 330062 365854
rect 330146 365618 330382 365854
rect 329826 365298 330062 365534
rect 330146 365298 330382 365534
rect 365826 365618 366062 365854
rect 366146 365618 366382 365854
rect 365826 365298 366062 365534
rect 366146 365298 366382 365534
rect 401826 365618 402062 365854
rect 402146 365618 402382 365854
rect 401826 365298 402062 365534
rect 402146 365298 402382 365534
rect 437826 365618 438062 365854
rect 438146 365618 438382 365854
rect 437826 365298 438062 365534
rect 438146 365298 438382 365534
rect 473826 365618 474062 365854
rect 474146 365618 474382 365854
rect 473826 365298 474062 365534
rect 474146 365298 474382 365534
rect 509826 365618 510062 365854
rect 510146 365618 510382 365854
rect 509826 365298 510062 365534
rect 510146 365298 510382 365534
rect 545826 365618 546062 365854
rect 546146 365618 546382 365854
rect 545826 365298 546062 365534
rect 546146 365298 546382 365534
rect 13198 334118 13434 334354
rect 13518 334118 13754 334354
rect 13198 333798 13434 334034
rect 13518 333798 13754 334034
rect 167826 334118 168062 334354
rect 168146 334118 168382 334354
rect 167826 333798 168062 334034
rect 168146 333798 168382 334034
rect 203826 334118 204062 334354
rect 204146 334118 204382 334354
rect 203826 333798 204062 334034
rect 204146 333798 204382 334034
rect 239826 334118 240062 334354
rect 240146 334118 240382 334354
rect 239826 333798 240062 334034
rect 240146 333798 240382 334034
rect 275826 334118 276062 334354
rect 276146 334118 276382 334354
rect 275826 333798 276062 334034
rect 276146 333798 276382 334034
rect 311826 334118 312062 334354
rect 312146 334118 312382 334354
rect 311826 333798 312062 334034
rect 312146 333798 312382 334034
rect 347826 334118 348062 334354
rect 348146 334118 348382 334354
rect 347826 333798 348062 334034
rect 348146 333798 348382 334034
rect 383826 334118 384062 334354
rect 384146 334118 384382 334354
rect 383826 333798 384062 334034
rect 384146 333798 384382 334034
rect 419826 334118 420062 334354
rect 420146 334118 420382 334354
rect 419826 333798 420062 334034
rect 420146 333798 420382 334034
rect 563826 334118 564062 334354
rect 564146 334118 564382 334354
rect 563826 333798 564062 334034
rect 564146 333798 564382 334034
rect 582326 334118 582562 334354
rect 582646 334118 582882 334354
rect 582326 333798 582562 334034
rect 582646 333798 582882 334034
rect -1974 329618 -1738 329854
rect -1654 329618 -1418 329854
rect -1974 329298 -1738 329534
rect -1654 329298 -1418 329534
rect 5826 329618 6062 329854
rect 6146 329618 6382 329854
rect 5826 329298 6062 329534
rect 6146 329298 6382 329534
rect 185826 329618 186062 329854
rect 186146 329618 186382 329854
rect 185826 329298 186062 329534
rect 186146 329298 186382 329534
rect 221826 329618 222062 329854
rect 222146 329618 222382 329854
rect 221826 329298 222062 329534
rect 222146 329298 222382 329534
rect 257826 329618 258062 329854
rect 258146 329618 258382 329854
rect 257826 329298 258062 329534
rect 258146 329298 258382 329534
rect 293826 329618 294062 329854
rect 294146 329618 294382 329854
rect 293826 329298 294062 329534
rect 294146 329298 294382 329534
rect 329826 329618 330062 329854
rect 330146 329618 330382 329854
rect 329826 329298 330062 329534
rect 330146 329298 330382 329534
rect 365826 329618 366062 329854
rect 366146 329618 366382 329854
rect 365826 329298 366062 329534
rect 366146 329298 366382 329534
rect 401826 329618 402062 329854
rect 402146 329618 402382 329854
rect 401826 329298 402062 329534
rect 402146 329298 402382 329534
rect 570350 329618 570586 329854
rect 570670 329618 570906 329854
rect 570350 329298 570586 329534
rect 570670 329298 570906 329534
rect 13198 298118 13434 298354
rect 13518 298118 13754 298354
rect 13198 297798 13434 298034
rect 13518 297798 13754 298034
rect 167826 298118 168062 298354
rect 168146 298118 168382 298354
rect 167826 297798 168062 298034
rect 168146 297798 168382 298034
rect 203826 298118 204062 298354
rect 204146 298118 204382 298354
rect 203826 297798 204062 298034
rect 204146 297798 204382 298034
rect 239826 298118 240062 298354
rect 240146 298118 240382 298354
rect 239826 297798 240062 298034
rect 240146 297798 240382 298034
rect 275826 298118 276062 298354
rect 276146 298118 276382 298354
rect 275826 297798 276062 298034
rect 276146 297798 276382 298034
rect 311826 298118 312062 298354
rect 312146 298118 312382 298354
rect 311826 297798 312062 298034
rect 312146 297798 312382 298034
rect 347826 298118 348062 298354
rect 348146 298118 348382 298354
rect 347826 297798 348062 298034
rect 348146 297798 348382 298034
rect 383826 298118 384062 298354
rect 384146 298118 384382 298354
rect 383826 297798 384062 298034
rect 384146 297798 384382 298034
rect 419826 298118 420062 298354
rect 420146 298118 420382 298354
rect 419826 297798 420062 298034
rect 420146 297798 420382 298034
rect 563826 298118 564062 298354
rect 564146 298118 564382 298354
rect 563826 297798 564062 298034
rect 564146 297798 564382 298034
rect 582326 298118 582562 298354
rect 582646 298118 582882 298354
rect 582326 297798 582562 298034
rect 582646 297798 582882 298034
rect -1974 293618 -1738 293854
rect -1654 293618 -1418 293854
rect -1974 293298 -1738 293534
rect -1654 293298 -1418 293534
rect 5826 293618 6062 293854
rect 6146 293618 6382 293854
rect 5826 293298 6062 293534
rect 6146 293298 6382 293534
rect 185826 293618 186062 293854
rect 186146 293618 186382 293854
rect 185826 293298 186062 293534
rect 186146 293298 186382 293534
rect 221826 293618 222062 293854
rect 222146 293618 222382 293854
rect 221826 293298 222062 293534
rect 222146 293298 222382 293534
rect 257826 293618 258062 293854
rect 258146 293618 258382 293854
rect 257826 293298 258062 293534
rect 258146 293298 258382 293534
rect 293826 293618 294062 293854
rect 294146 293618 294382 293854
rect 293826 293298 294062 293534
rect 294146 293298 294382 293534
rect 329826 293618 330062 293854
rect 330146 293618 330382 293854
rect 329826 293298 330062 293534
rect 330146 293298 330382 293534
rect 365826 293618 366062 293854
rect 366146 293618 366382 293854
rect 365826 293298 366062 293534
rect 366146 293298 366382 293534
rect 401826 293618 402062 293854
rect 402146 293618 402382 293854
rect 401826 293298 402062 293534
rect 402146 293298 402382 293534
rect 570350 293618 570586 293854
rect 570670 293618 570906 293854
rect 570350 293298 570586 293534
rect 570670 293298 570906 293534
rect 13198 262118 13434 262354
rect 13518 262118 13754 262354
rect 13198 261798 13434 262034
rect 13518 261798 13754 262034
rect 167826 262118 168062 262354
rect 168146 262118 168382 262354
rect 167826 261798 168062 262034
rect 168146 261798 168382 262034
rect 203826 262118 204062 262354
rect 204146 262118 204382 262354
rect 203826 261798 204062 262034
rect 204146 261798 204382 262034
rect 239826 262118 240062 262354
rect 240146 262118 240382 262354
rect 239826 261798 240062 262034
rect 240146 261798 240382 262034
rect 275826 262118 276062 262354
rect 276146 262118 276382 262354
rect 275826 261798 276062 262034
rect 276146 261798 276382 262034
rect 311826 262118 312062 262354
rect 312146 262118 312382 262354
rect 311826 261798 312062 262034
rect 312146 261798 312382 262034
rect 347826 262118 348062 262354
rect 348146 262118 348382 262354
rect 347826 261798 348062 262034
rect 348146 261798 348382 262034
rect 383826 262118 384062 262354
rect 384146 262118 384382 262354
rect 383826 261798 384062 262034
rect 384146 261798 384382 262034
rect 419826 262118 420062 262354
rect 420146 262118 420382 262354
rect 419826 261798 420062 262034
rect 420146 261798 420382 262034
rect 563826 262118 564062 262354
rect 564146 262118 564382 262354
rect 563826 261798 564062 262034
rect 564146 261798 564382 262034
rect 582326 262118 582562 262354
rect 582646 262118 582882 262354
rect 582326 261798 582562 262034
rect 582646 261798 582882 262034
rect -1974 257618 -1738 257854
rect -1654 257618 -1418 257854
rect -1974 257298 -1738 257534
rect -1654 257298 -1418 257534
rect 5826 257618 6062 257854
rect 6146 257618 6382 257854
rect 5826 257298 6062 257534
rect 6146 257298 6382 257534
rect 185826 257618 186062 257854
rect 186146 257618 186382 257854
rect 185826 257298 186062 257534
rect 186146 257298 186382 257534
rect 221826 257618 222062 257854
rect 222146 257618 222382 257854
rect 221826 257298 222062 257534
rect 222146 257298 222382 257534
rect 257826 257618 258062 257854
rect 258146 257618 258382 257854
rect 257826 257298 258062 257534
rect 258146 257298 258382 257534
rect 293826 257618 294062 257854
rect 294146 257618 294382 257854
rect 293826 257298 294062 257534
rect 294146 257298 294382 257534
rect 329826 257618 330062 257854
rect 330146 257618 330382 257854
rect 329826 257298 330062 257534
rect 330146 257298 330382 257534
rect 365826 257618 366062 257854
rect 366146 257618 366382 257854
rect 365826 257298 366062 257534
rect 366146 257298 366382 257534
rect 401826 257618 402062 257854
rect 402146 257618 402382 257854
rect 401826 257298 402062 257534
rect 402146 257298 402382 257534
rect 570350 257618 570586 257854
rect 570670 257618 570906 257854
rect 570350 257298 570586 257534
rect 570670 257298 570906 257534
rect 23826 226118 24062 226354
rect 24146 226118 24382 226354
rect 23826 225798 24062 226034
rect 24146 225798 24382 226034
rect 59826 226118 60062 226354
rect 60146 226118 60382 226354
rect 59826 225798 60062 226034
rect 60146 225798 60382 226034
rect 95826 226118 96062 226354
rect 96146 226118 96382 226354
rect 95826 225798 96062 226034
rect 96146 225798 96382 226034
rect 131826 226118 132062 226354
rect 132146 226118 132382 226354
rect 131826 225798 132062 226034
rect 132146 225798 132382 226034
rect 167826 226118 168062 226354
rect 168146 226118 168382 226354
rect 167826 225798 168062 226034
rect 168146 225798 168382 226034
rect 203826 226118 204062 226354
rect 204146 226118 204382 226354
rect 203826 225798 204062 226034
rect 204146 225798 204382 226034
rect 239826 226118 240062 226354
rect 240146 226118 240382 226354
rect 239826 225798 240062 226034
rect 240146 225798 240382 226034
rect 275826 226118 276062 226354
rect 276146 226118 276382 226354
rect 275826 225798 276062 226034
rect 276146 225798 276382 226034
rect 311826 226118 312062 226354
rect 312146 226118 312382 226354
rect 311826 225798 312062 226034
rect 312146 225798 312382 226034
rect 347826 226118 348062 226354
rect 348146 226118 348382 226354
rect 347826 225798 348062 226034
rect 348146 225798 348382 226034
rect 383826 226118 384062 226354
rect 384146 226118 384382 226354
rect 383826 225798 384062 226034
rect 384146 225798 384382 226034
rect 419826 226118 420062 226354
rect 420146 226118 420382 226354
rect 419826 225798 420062 226034
rect 420146 225798 420382 226034
rect 455826 226118 456062 226354
rect 456146 226118 456382 226354
rect 455826 225798 456062 226034
rect 456146 225798 456382 226034
rect 491826 226118 492062 226354
rect 492146 226118 492382 226354
rect 491826 225798 492062 226034
rect 492146 225798 492382 226034
rect 527826 226118 528062 226354
rect 528146 226118 528382 226354
rect 527826 225798 528062 226034
rect 528146 225798 528382 226034
rect 563826 226118 564062 226354
rect 564146 226118 564382 226354
rect 563826 225798 564062 226034
rect 564146 225798 564382 226034
rect 582326 226118 582562 226354
rect 582646 226118 582882 226354
rect 582326 225798 582562 226034
rect 582646 225798 582882 226034
rect -1974 221618 -1738 221854
rect -1654 221618 -1418 221854
rect -1974 221298 -1738 221534
rect -1654 221298 -1418 221534
rect 5826 221618 6062 221854
rect 6146 221618 6382 221854
rect 5826 221298 6062 221534
rect 6146 221298 6382 221534
rect 185826 221618 186062 221854
rect 186146 221618 186382 221854
rect 185826 221298 186062 221534
rect 186146 221298 186382 221534
rect 221826 221618 222062 221854
rect 222146 221618 222382 221854
rect 221826 221298 222062 221534
rect 222146 221298 222382 221534
rect 257826 221618 258062 221854
rect 258146 221618 258382 221854
rect 257826 221298 258062 221534
rect 258146 221298 258382 221534
rect 293826 221618 294062 221854
rect 294146 221618 294382 221854
rect 293826 221298 294062 221534
rect 294146 221298 294382 221534
rect 329826 221618 330062 221854
rect 330146 221618 330382 221854
rect 329826 221298 330062 221534
rect 330146 221298 330382 221534
rect 365826 221618 366062 221854
rect 366146 221618 366382 221854
rect 365826 221298 366062 221534
rect 366146 221298 366382 221534
rect 401826 221618 402062 221854
rect 402146 221618 402382 221854
rect 401826 221298 402062 221534
rect 402146 221298 402382 221534
rect 570350 221618 570586 221854
rect 570670 221618 570906 221854
rect 570350 221298 570586 221534
rect 570670 221298 570906 221534
rect 13198 190118 13434 190354
rect 13518 190118 13754 190354
rect 13198 189798 13434 190034
rect 13518 189798 13754 190034
rect 167826 190118 168062 190354
rect 168146 190118 168382 190354
rect 167826 189798 168062 190034
rect 168146 189798 168382 190034
rect 203826 190118 204062 190354
rect 204146 190118 204382 190354
rect 203826 189798 204062 190034
rect 204146 189798 204382 190034
rect 239826 190118 240062 190354
rect 240146 190118 240382 190354
rect 239826 189798 240062 190034
rect 240146 189798 240382 190034
rect 275826 190118 276062 190354
rect 276146 190118 276382 190354
rect 275826 189798 276062 190034
rect 276146 189798 276382 190034
rect 311826 190118 312062 190354
rect 312146 190118 312382 190354
rect 311826 189798 312062 190034
rect 312146 189798 312382 190034
rect 347826 190118 348062 190354
rect 348146 190118 348382 190354
rect 347826 189798 348062 190034
rect 348146 189798 348382 190034
rect 383826 190118 384062 190354
rect 384146 190118 384382 190354
rect 383826 189798 384062 190034
rect 384146 189798 384382 190034
rect 419826 190118 420062 190354
rect 420146 190118 420382 190354
rect 419826 189798 420062 190034
rect 420146 189798 420382 190034
rect 563826 190118 564062 190354
rect 564146 190118 564382 190354
rect 563826 189798 564062 190034
rect 564146 189798 564382 190034
rect 582326 190118 582562 190354
rect 582646 190118 582882 190354
rect 582326 189798 582562 190034
rect 582646 189798 582882 190034
rect -1974 185618 -1738 185854
rect -1654 185618 -1418 185854
rect -1974 185298 -1738 185534
rect -1654 185298 -1418 185534
rect 5826 185618 6062 185854
rect 6146 185618 6382 185854
rect 5826 185298 6062 185534
rect 6146 185298 6382 185534
rect 185826 185618 186062 185854
rect 186146 185618 186382 185854
rect 185826 185298 186062 185534
rect 186146 185298 186382 185534
rect 221826 185618 222062 185854
rect 222146 185618 222382 185854
rect 221826 185298 222062 185534
rect 222146 185298 222382 185534
rect 257826 185618 258062 185854
rect 258146 185618 258382 185854
rect 257826 185298 258062 185534
rect 258146 185298 258382 185534
rect 293826 185618 294062 185854
rect 294146 185618 294382 185854
rect 293826 185298 294062 185534
rect 294146 185298 294382 185534
rect 329826 185618 330062 185854
rect 330146 185618 330382 185854
rect 329826 185298 330062 185534
rect 330146 185298 330382 185534
rect 365826 185618 366062 185854
rect 366146 185618 366382 185854
rect 365826 185298 366062 185534
rect 366146 185298 366382 185534
rect 401826 185618 402062 185854
rect 402146 185618 402382 185854
rect 401826 185298 402062 185534
rect 402146 185298 402382 185534
rect 570350 185618 570586 185854
rect 570670 185618 570906 185854
rect 570350 185298 570586 185534
rect 570670 185298 570906 185534
rect 13198 154118 13434 154354
rect 13518 154118 13754 154354
rect 13198 153798 13434 154034
rect 13518 153798 13754 154034
rect 167826 154118 168062 154354
rect 168146 154118 168382 154354
rect 167826 153798 168062 154034
rect 168146 153798 168382 154034
rect 203826 154118 204062 154354
rect 204146 154118 204382 154354
rect 203826 153798 204062 154034
rect 204146 153798 204382 154034
rect 239826 154118 240062 154354
rect 240146 154118 240382 154354
rect 239826 153798 240062 154034
rect 240146 153798 240382 154034
rect 275826 154118 276062 154354
rect 276146 154118 276382 154354
rect 275826 153798 276062 154034
rect 276146 153798 276382 154034
rect 311826 154118 312062 154354
rect 312146 154118 312382 154354
rect 311826 153798 312062 154034
rect 312146 153798 312382 154034
rect 347826 154118 348062 154354
rect 348146 154118 348382 154354
rect 347826 153798 348062 154034
rect 348146 153798 348382 154034
rect 383826 154118 384062 154354
rect 384146 154118 384382 154354
rect 383826 153798 384062 154034
rect 384146 153798 384382 154034
rect 419826 154118 420062 154354
rect 420146 154118 420382 154354
rect 419826 153798 420062 154034
rect 420146 153798 420382 154034
rect 563826 154118 564062 154354
rect 564146 154118 564382 154354
rect 563826 153798 564062 154034
rect 564146 153798 564382 154034
rect 582326 154118 582562 154354
rect 582646 154118 582882 154354
rect 582326 153798 582562 154034
rect 582646 153798 582882 154034
rect -1974 149618 -1738 149854
rect -1654 149618 -1418 149854
rect -1974 149298 -1738 149534
rect -1654 149298 -1418 149534
rect 5826 149618 6062 149854
rect 6146 149618 6382 149854
rect 5826 149298 6062 149534
rect 6146 149298 6382 149534
rect 185826 149618 186062 149854
rect 186146 149618 186382 149854
rect 185826 149298 186062 149534
rect 186146 149298 186382 149534
rect 221826 149618 222062 149854
rect 222146 149618 222382 149854
rect 221826 149298 222062 149534
rect 222146 149298 222382 149534
rect 257826 149618 258062 149854
rect 258146 149618 258382 149854
rect 257826 149298 258062 149534
rect 258146 149298 258382 149534
rect 293826 149618 294062 149854
rect 294146 149618 294382 149854
rect 293826 149298 294062 149534
rect 294146 149298 294382 149534
rect 329826 149618 330062 149854
rect 330146 149618 330382 149854
rect 329826 149298 330062 149534
rect 330146 149298 330382 149534
rect 365826 149618 366062 149854
rect 366146 149618 366382 149854
rect 365826 149298 366062 149534
rect 366146 149298 366382 149534
rect 401826 149618 402062 149854
rect 402146 149618 402382 149854
rect 401826 149298 402062 149534
rect 402146 149298 402382 149534
rect 570350 149618 570586 149854
rect 570670 149618 570906 149854
rect 570350 149298 570586 149534
rect 570670 149298 570906 149534
rect 23826 118118 24062 118354
rect 24146 118118 24382 118354
rect 23826 117798 24062 118034
rect 24146 117798 24382 118034
rect 59826 118118 60062 118354
rect 60146 118118 60382 118354
rect 59826 117798 60062 118034
rect 60146 117798 60382 118034
rect 95826 118118 96062 118354
rect 96146 118118 96382 118354
rect 95826 117798 96062 118034
rect 96146 117798 96382 118034
rect 131826 118118 132062 118354
rect 132146 118118 132382 118354
rect 131826 117798 132062 118034
rect 132146 117798 132382 118034
rect 167826 118118 168062 118354
rect 168146 118118 168382 118354
rect 167826 117798 168062 118034
rect 168146 117798 168382 118034
rect 203826 118118 204062 118354
rect 204146 118118 204382 118354
rect 203826 117798 204062 118034
rect 204146 117798 204382 118034
rect 239826 118118 240062 118354
rect 240146 118118 240382 118354
rect 239826 117798 240062 118034
rect 240146 117798 240382 118034
rect 275826 118118 276062 118354
rect 276146 118118 276382 118354
rect 275826 117798 276062 118034
rect 276146 117798 276382 118034
rect 311826 118118 312062 118354
rect 312146 118118 312382 118354
rect 311826 117798 312062 118034
rect 312146 117798 312382 118034
rect 347826 118118 348062 118354
rect 348146 118118 348382 118354
rect 347826 117798 348062 118034
rect 348146 117798 348382 118034
rect 383826 118118 384062 118354
rect 384146 118118 384382 118354
rect 383826 117798 384062 118034
rect 384146 117798 384382 118034
rect 419826 118118 420062 118354
rect 420146 118118 420382 118354
rect 419826 117798 420062 118034
rect 420146 117798 420382 118034
rect 455826 118118 456062 118354
rect 456146 118118 456382 118354
rect 455826 117798 456062 118034
rect 456146 117798 456382 118034
rect 491826 118118 492062 118354
rect 492146 118118 492382 118354
rect 491826 117798 492062 118034
rect 492146 117798 492382 118034
rect 527826 118118 528062 118354
rect 528146 118118 528382 118354
rect 527826 117798 528062 118034
rect 528146 117798 528382 118034
rect 563826 118118 564062 118354
rect 564146 118118 564382 118354
rect 563826 117798 564062 118034
rect 564146 117798 564382 118034
rect 582326 118118 582562 118354
rect 582646 118118 582882 118354
rect 582326 117798 582562 118034
rect 582646 117798 582882 118034
rect -1974 113618 -1738 113854
rect -1654 113618 -1418 113854
rect -1974 113298 -1738 113534
rect -1654 113298 -1418 113534
rect 5826 113618 6062 113854
rect 6146 113618 6382 113854
rect 5826 113298 6062 113534
rect 6146 113298 6382 113534
rect 41826 113479 42062 113715
rect 42146 113479 42382 113715
rect 77826 113479 78062 113715
rect 78146 113479 78382 113715
rect 113826 113479 114062 113715
rect 114146 113479 114382 113715
rect 149826 113479 150062 113715
rect 150146 113479 150382 113715
rect 293826 113618 294062 113854
rect 294146 113618 294382 113854
rect 293826 113298 294062 113534
rect 294146 113298 294382 113534
rect 401826 113618 402062 113854
rect 402146 113618 402382 113854
rect 401826 113298 402062 113534
rect 402146 113298 402382 113534
rect 437826 113479 438062 113715
rect 438146 113479 438382 113715
rect 473826 113479 474062 113715
rect 474146 113479 474382 113715
rect 509826 113479 510062 113715
rect 510146 113479 510382 113715
rect 545826 113479 546062 113715
rect 546146 113479 546382 113715
rect 13198 82118 13434 82354
rect 13518 82118 13754 82354
rect 13198 81798 13434 82034
rect 13518 81798 13754 82034
rect 167826 82118 168062 82354
rect 168146 82118 168382 82354
rect 167826 81798 168062 82034
rect 168146 81798 168382 82034
rect 291590 82118 291826 82354
rect 291910 82118 292146 82354
rect 291590 81798 291826 82034
rect 291910 81798 292146 82034
rect 419826 82118 420062 82354
rect 420146 82118 420382 82354
rect 419826 81798 420062 82034
rect 420146 81798 420382 82034
rect 563826 82118 564062 82354
rect 564146 82118 564382 82354
rect 563826 81798 564062 82034
rect 564146 81798 564382 82034
rect 582326 82118 582562 82354
rect 582646 82118 582882 82354
rect 582326 81798 582562 82034
rect 582646 81798 582882 82034
rect -1974 77618 -1738 77854
rect -1654 77618 -1418 77854
rect -1974 77298 -1738 77534
rect -1654 77298 -1418 77534
rect 5826 77618 6062 77854
rect 6146 77618 6382 77854
rect 5826 77298 6062 77534
rect 6146 77298 6382 77534
rect 173094 77618 173330 77854
rect 173414 77618 173650 77854
rect 173094 77298 173330 77534
rect 173414 77298 173650 77534
rect 293826 77618 294062 77854
rect 294146 77618 294382 77854
rect 293826 77298 294062 77534
rect 294146 77298 294382 77534
rect 401826 77618 402062 77854
rect 402146 77618 402382 77854
rect 401826 77298 402062 77534
rect 402146 77298 402382 77534
rect 570350 77618 570586 77854
rect 570670 77618 570906 77854
rect 570350 77298 570586 77534
rect 570670 77298 570906 77534
rect 13198 46118 13434 46354
rect 13518 46118 13754 46354
rect 13198 45798 13434 46034
rect 13518 45798 13754 46034
rect 167826 46118 168062 46354
rect 168146 46118 168382 46354
rect 167826 45798 168062 46034
rect 168146 45798 168382 46034
rect 291590 46118 291826 46354
rect 291910 46118 292146 46354
rect 291590 45798 291826 46034
rect 291910 45798 292146 46034
rect 419826 46118 420062 46354
rect 420146 46118 420382 46354
rect 419826 45798 420062 46034
rect 420146 45798 420382 46034
rect 563826 46118 564062 46354
rect 564146 46118 564382 46354
rect 563826 45798 564062 46034
rect 564146 45798 564382 46034
rect 582326 46118 582562 46354
rect 582646 46118 582882 46354
rect 582326 45798 582562 46034
rect 582646 45798 582882 46034
rect -1974 41618 -1738 41854
rect -1654 41618 -1418 41854
rect -1974 41298 -1738 41534
rect -1654 41298 -1418 41534
rect 5826 41618 6062 41854
rect 6146 41618 6382 41854
rect 5826 41298 6062 41534
rect 6146 41298 6382 41534
rect 173094 41618 173330 41854
rect 173414 41618 173650 41854
rect 173094 41298 173330 41534
rect 173414 41298 173650 41534
rect 293826 41618 294062 41854
rect 294146 41618 294382 41854
rect 293826 41298 294062 41534
rect 294146 41298 294382 41534
rect 401826 41618 402062 41854
rect 402146 41618 402382 41854
rect 401826 41298 402062 41534
rect 402146 41298 402382 41534
rect 570350 41618 570586 41854
rect 570670 41618 570906 41854
rect 570350 41298 570586 41534
rect 570670 41298 570906 41534
rect 23826 10118 24062 10354
rect 24146 10118 24382 10354
rect 23826 9798 24062 10034
rect 24146 9798 24382 10034
rect 59826 10118 60062 10354
rect 60146 10118 60382 10354
rect 59826 9798 60062 10034
rect 60146 9798 60382 10034
rect 95826 10118 96062 10354
rect 96146 10118 96382 10354
rect 95826 9798 96062 10034
rect 96146 9798 96382 10034
rect 131826 10118 132062 10354
rect 132146 10118 132382 10354
rect 131826 9798 132062 10034
rect 132146 9798 132382 10034
rect 167826 10118 168062 10354
rect 168146 10118 168382 10354
rect 167826 9798 168062 10034
rect 168146 9798 168382 10034
rect 203826 10118 204062 10354
rect 204146 10118 204382 10354
rect 203826 9798 204062 10034
rect 204146 9798 204382 10034
rect 239826 10118 240062 10354
rect 240146 10118 240382 10354
rect 239826 9798 240062 10034
rect 240146 9798 240382 10034
rect 275826 10118 276062 10354
rect 276146 10118 276382 10354
rect 275826 9798 276062 10034
rect 276146 9798 276382 10034
rect 311826 10118 312062 10354
rect 312146 10118 312382 10354
rect 311826 9798 312062 10034
rect 312146 9798 312382 10034
rect 347826 10118 348062 10354
rect 348146 10118 348382 10354
rect 347826 9798 348062 10034
rect 348146 9798 348382 10034
rect 383826 10118 384062 10354
rect 384146 10118 384382 10354
rect 383826 9798 384062 10034
rect 384146 9798 384382 10034
rect 419826 10118 420062 10354
rect 420146 10118 420382 10354
rect 419826 9798 420062 10034
rect 420146 9798 420382 10034
rect 455826 10118 456062 10354
rect 456146 10118 456382 10354
rect 455826 9798 456062 10034
rect 456146 9798 456382 10034
rect 491826 10118 492062 10354
rect 492146 10118 492382 10354
rect 491826 9798 492062 10034
rect 492146 9798 492382 10034
rect 527826 10118 528062 10354
rect 528146 10118 528382 10354
rect 527826 9798 528062 10034
rect 528146 9798 528382 10034
rect 563826 10118 564062 10354
rect 564146 10118 564382 10354
rect 563826 9798 564062 10034
rect 564146 9798 564382 10034
rect 582326 10118 582562 10354
rect 582646 10118 582882 10354
rect 582326 9798 582562 10034
rect 582646 9798 582882 10034
rect -1974 5618 -1738 5854
rect -1654 5618 -1418 5854
rect -1974 5298 -1738 5534
rect -1654 5298 -1418 5534
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 689618 585578 689854
rect 585662 689618 585898 689854
rect 585342 689298 585578 689534
rect 585662 689298 585898 689534
rect 585342 653618 585578 653854
rect 585662 653618 585898 653854
rect 585342 653298 585578 653534
rect 585662 653298 585898 653534
rect 585342 617618 585578 617854
rect 585662 617618 585898 617854
rect 585342 617298 585578 617534
rect 585662 617298 585898 617534
rect 585342 581618 585578 581854
rect 585662 581618 585898 581854
rect 585342 581298 585578 581534
rect 585662 581298 585898 581534
rect 585342 545618 585578 545854
rect 585662 545618 585898 545854
rect 585342 545298 585578 545534
rect 585662 545298 585898 545534
rect 585342 509618 585578 509854
rect 585662 509618 585898 509854
rect 585342 509298 585578 509534
rect 585662 509298 585898 509534
rect 585342 473618 585578 473854
rect 585662 473618 585898 473854
rect 585342 473298 585578 473534
rect 585662 473298 585898 473534
rect 585342 437618 585578 437854
rect 585662 437618 585898 437854
rect 585342 437298 585578 437534
rect 585662 437298 585898 437534
rect 585342 401618 585578 401854
rect 585662 401618 585898 401854
rect 585342 401298 585578 401534
rect 585662 401298 585898 401534
rect 585342 365618 585578 365854
rect 585662 365618 585898 365854
rect 585342 365298 585578 365534
rect 585662 365298 585898 365534
rect 585342 329618 585578 329854
rect 585662 329618 585898 329854
rect 585342 329298 585578 329534
rect 585662 329298 585898 329534
rect 585342 293618 585578 293854
rect 585662 293618 585898 293854
rect 585342 293298 585578 293534
rect 585662 293298 585898 293534
rect 585342 257618 585578 257854
rect 585662 257618 585898 257854
rect 585342 257298 585578 257534
rect 585662 257298 585898 257534
rect 585342 221618 585578 221854
rect 585662 221618 585898 221854
rect 585342 221298 585578 221534
rect 585662 221298 585898 221534
rect 585342 185618 585578 185854
rect 585662 185618 585898 185854
rect 585342 185298 585578 185534
rect 585662 185298 585898 185534
rect 585342 149618 585578 149854
rect 585662 149618 585898 149854
rect 585342 149298 585578 149534
rect 585662 149298 585898 149534
rect 585342 113618 585578 113854
rect 585662 113618 585898 113854
rect 585342 113298 585578 113534
rect 585662 113298 585898 113534
rect 585342 77618 585578 77854
rect 585662 77618 585898 77854
rect 585342 77298 585578 77534
rect 585662 77298 585898 77534
rect 585342 41618 585578 41854
rect 585662 41618 585898 41854
rect 585342 41298 585578 41534
rect 585662 41298 585898 41534
rect 585342 5618 585578 5854
rect 585662 5618 585898 5854
rect 585342 5298 585578 5534
rect 585662 5298 585898 5534
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 694118 586538 694354
rect 586622 694118 586858 694354
rect 586302 693798 586538 694034
rect 586622 693798 586858 694034
rect 586302 658118 586538 658354
rect 586622 658118 586858 658354
rect 586302 657798 586538 658034
rect 586622 657798 586858 658034
rect 586302 622118 586538 622354
rect 586622 622118 586858 622354
rect 586302 621798 586538 622034
rect 586622 621798 586858 622034
rect 586302 586118 586538 586354
rect 586622 586118 586858 586354
rect 586302 585798 586538 586034
rect 586622 585798 586858 586034
rect 586302 550118 586538 550354
rect 586622 550118 586858 550354
rect 586302 549798 586538 550034
rect 586622 549798 586858 550034
rect 586302 514118 586538 514354
rect 586622 514118 586858 514354
rect 586302 513798 586538 514034
rect 586622 513798 586858 514034
rect 586302 478118 586538 478354
rect 586622 478118 586858 478354
rect 586302 477798 586538 478034
rect 586622 477798 586858 478034
rect 586302 442118 586538 442354
rect 586622 442118 586858 442354
rect 586302 441798 586538 442034
rect 586622 441798 586858 442034
rect 586302 406118 586538 406354
rect 586622 406118 586858 406354
rect 586302 405798 586538 406034
rect 586622 405798 586858 406034
rect 586302 370118 586538 370354
rect 586622 370118 586858 370354
rect 586302 369798 586538 370034
rect 586622 369798 586858 370034
rect 586302 334118 586538 334354
rect 586622 334118 586858 334354
rect 586302 333798 586538 334034
rect 586622 333798 586858 334034
rect 586302 298118 586538 298354
rect 586622 298118 586858 298354
rect 586302 297798 586538 298034
rect 586622 297798 586858 298034
rect 586302 262118 586538 262354
rect 586622 262118 586858 262354
rect 586302 261798 586538 262034
rect 586622 261798 586858 262034
rect 586302 226118 586538 226354
rect 586622 226118 586858 226354
rect 586302 225798 586538 226034
rect 586622 225798 586858 226034
rect 586302 190118 586538 190354
rect 586622 190118 586858 190354
rect 586302 189798 586538 190034
rect 586622 189798 586858 190034
rect 586302 154118 586538 154354
rect 586622 154118 586858 154354
rect 586302 153798 586538 154034
rect 586622 153798 586858 154034
rect 586302 118118 586538 118354
rect 586622 118118 586858 118354
rect 586302 117798 586538 118034
rect 586622 117798 586858 118034
rect 586302 82118 586538 82354
rect 586622 82118 586858 82354
rect 586302 81798 586538 82034
rect 586622 81798 586858 82034
rect 586302 46118 586538 46354
rect 586622 46118 586858 46354
rect 586302 45798 586538 46034
rect 586622 45798 586858 46034
rect 586302 10118 586538 10354
rect 586622 10118 586858 10354
rect 586302 9798 586538 10034
rect 586622 9798 586858 10034
rect 582326 -1542 582562 -1306
rect 582646 -1542 582882 -1306
rect 582326 -1862 582562 -1626
rect 582646 -1862 582882 -1626
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 582326 705798
rect 582562 705562 582646 705798
rect 582882 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 582326 705478
rect 582562 705242 582646 705478
rect 582882 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 694354 592650 694386
rect -8726 694118 -2934 694354
rect -2698 694118 -2614 694354
rect -2378 694118 23826 694354
rect 24062 694118 24146 694354
rect 24382 694118 59826 694354
rect 60062 694118 60146 694354
rect 60382 694118 95826 694354
rect 96062 694118 96146 694354
rect 96382 694118 131826 694354
rect 132062 694118 132146 694354
rect 132382 694118 167826 694354
rect 168062 694118 168146 694354
rect 168382 694118 203826 694354
rect 204062 694118 204146 694354
rect 204382 694118 239826 694354
rect 240062 694118 240146 694354
rect 240382 694118 275826 694354
rect 276062 694118 276146 694354
rect 276382 694118 311826 694354
rect 312062 694118 312146 694354
rect 312382 694118 347826 694354
rect 348062 694118 348146 694354
rect 348382 694118 383826 694354
rect 384062 694118 384146 694354
rect 384382 694118 419826 694354
rect 420062 694118 420146 694354
rect 420382 694118 455826 694354
rect 456062 694118 456146 694354
rect 456382 694118 491826 694354
rect 492062 694118 492146 694354
rect 492382 694118 527826 694354
rect 528062 694118 528146 694354
rect 528382 694118 563826 694354
rect 564062 694118 564146 694354
rect 564382 694118 582326 694354
rect 582562 694118 582646 694354
rect 582882 694118 586302 694354
rect 586538 694118 586622 694354
rect 586858 694118 592650 694354
rect -8726 694034 592650 694118
rect -8726 693798 -2934 694034
rect -2698 693798 -2614 694034
rect -2378 693798 23826 694034
rect 24062 693798 24146 694034
rect 24382 693798 59826 694034
rect 60062 693798 60146 694034
rect 60382 693798 95826 694034
rect 96062 693798 96146 694034
rect 96382 693798 131826 694034
rect 132062 693798 132146 694034
rect 132382 693798 167826 694034
rect 168062 693798 168146 694034
rect 168382 693798 203826 694034
rect 204062 693798 204146 694034
rect 204382 693798 239826 694034
rect 240062 693798 240146 694034
rect 240382 693798 275826 694034
rect 276062 693798 276146 694034
rect 276382 693798 311826 694034
rect 312062 693798 312146 694034
rect 312382 693798 347826 694034
rect 348062 693798 348146 694034
rect 348382 693798 383826 694034
rect 384062 693798 384146 694034
rect 384382 693798 419826 694034
rect 420062 693798 420146 694034
rect 420382 693798 455826 694034
rect 456062 693798 456146 694034
rect 456382 693798 491826 694034
rect 492062 693798 492146 694034
rect 492382 693798 527826 694034
rect 528062 693798 528146 694034
rect 528382 693798 563826 694034
rect 564062 693798 564146 694034
rect 564382 693798 582326 694034
rect 582562 693798 582646 694034
rect 582882 693798 586302 694034
rect 586538 693798 586622 694034
rect 586858 693798 592650 694034
rect -8726 693766 592650 693798
rect -8726 689854 592650 689886
rect -8726 689618 -1974 689854
rect -1738 689618 -1654 689854
rect -1418 689618 5826 689854
rect 6062 689618 6146 689854
rect 6382 689618 41826 689854
rect 42062 689618 42146 689854
rect 42382 689618 77826 689854
rect 78062 689618 78146 689854
rect 78382 689618 113826 689854
rect 114062 689618 114146 689854
rect 114382 689618 149826 689854
rect 150062 689618 150146 689854
rect 150382 689618 185826 689854
rect 186062 689618 186146 689854
rect 186382 689618 221826 689854
rect 222062 689618 222146 689854
rect 222382 689618 257826 689854
rect 258062 689618 258146 689854
rect 258382 689618 293826 689854
rect 294062 689618 294146 689854
rect 294382 689618 329826 689854
rect 330062 689618 330146 689854
rect 330382 689618 365826 689854
rect 366062 689618 366146 689854
rect 366382 689618 401826 689854
rect 402062 689618 402146 689854
rect 402382 689618 437826 689854
rect 438062 689618 438146 689854
rect 438382 689618 473826 689854
rect 474062 689618 474146 689854
rect 474382 689618 509826 689854
rect 510062 689618 510146 689854
rect 510382 689618 545826 689854
rect 546062 689618 546146 689854
rect 546382 689618 585342 689854
rect 585578 689618 585662 689854
rect 585898 689618 592650 689854
rect -8726 689534 592650 689618
rect -8726 689298 -1974 689534
rect -1738 689298 -1654 689534
rect -1418 689298 5826 689534
rect 6062 689298 6146 689534
rect 6382 689298 41826 689534
rect 42062 689298 42146 689534
rect 42382 689298 77826 689534
rect 78062 689298 78146 689534
rect 78382 689298 113826 689534
rect 114062 689298 114146 689534
rect 114382 689298 149826 689534
rect 150062 689298 150146 689534
rect 150382 689298 185826 689534
rect 186062 689298 186146 689534
rect 186382 689298 221826 689534
rect 222062 689298 222146 689534
rect 222382 689298 257826 689534
rect 258062 689298 258146 689534
rect 258382 689298 293826 689534
rect 294062 689298 294146 689534
rect 294382 689298 329826 689534
rect 330062 689298 330146 689534
rect 330382 689298 365826 689534
rect 366062 689298 366146 689534
rect 366382 689298 401826 689534
rect 402062 689298 402146 689534
rect 402382 689298 437826 689534
rect 438062 689298 438146 689534
rect 438382 689298 473826 689534
rect 474062 689298 474146 689534
rect 474382 689298 509826 689534
rect 510062 689298 510146 689534
rect 510382 689298 545826 689534
rect 546062 689298 546146 689534
rect 546382 689298 585342 689534
rect 585578 689298 585662 689534
rect 585898 689298 592650 689534
rect -8726 689266 592650 689298
rect -8726 658354 592650 658386
rect -8726 658118 -2934 658354
rect -2698 658118 -2614 658354
rect -2378 658118 13198 658354
rect 13434 658118 13518 658354
rect 13754 658118 167826 658354
rect 168062 658118 168146 658354
rect 168382 658118 291590 658354
rect 291826 658118 291910 658354
rect 292146 658118 419826 658354
rect 420062 658118 420146 658354
rect 420382 658118 563826 658354
rect 564062 658118 564146 658354
rect 564382 658118 582326 658354
rect 582562 658118 582646 658354
rect 582882 658118 586302 658354
rect 586538 658118 586622 658354
rect 586858 658118 592650 658354
rect -8726 658034 592650 658118
rect -8726 657798 -2934 658034
rect -2698 657798 -2614 658034
rect -2378 657798 13198 658034
rect 13434 657798 13518 658034
rect 13754 657798 167826 658034
rect 168062 657798 168146 658034
rect 168382 657798 291590 658034
rect 291826 657798 291910 658034
rect 292146 657798 419826 658034
rect 420062 657798 420146 658034
rect 420382 657798 563826 658034
rect 564062 657798 564146 658034
rect 564382 657798 582326 658034
rect 582562 657798 582646 658034
rect 582882 657798 586302 658034
rect 586538 657798 586622 658034
rect 586858 657798 592650 658034
rect -8726 657766 592650 657798
rect -8726 653854 592650 653886
rect -8726 653618 -1974 653854
rect -1738 653618 -1654 653854
rect -1418 653618 5826 653854
rect 6062 653618 6146 653854
rect 6382 653618 173094 653854
rect 173330 653618 173414 653854
rect 173650 653618 293826 653854
rect 294062 653618 294146 653854
rect 294382 653618 401826 653854
rect 402062 653618 402146 653854
rect 402382 653618 570350 653854
rect 570586 653618 570670 653854
rect 570906 653618 585342 653854
rect 585578 653618 585662 653854
rect 585898 653618 592650 653854
rect -8726 653534 592650 653618
rect -8726 653298 -1974 653534
rect -1738 653298 -1654 653534
rect -1418 653298 5826 653534
rect 6062 653298 6146 653534
rect 6382 653298 173094 653534
rect 173330 653298 173414 653534
rect 173650 653298 293826 653534
rect 294062 653298 294146 653534
rect 294382 653298 401826 653534
rect 402062 653298 402146 653534
rect 402382 653298 570350 653534
rect 570586 653298 570670 653534
rect 570906 653298 585342 653534
rect 585578 653298 585662 653534
rect 585898 653298 592650 653534
rect -8726 653266 592650 653298
rect -8726 622354 592650 622386
rect -8726 622118 -2934 622354
rect -2698 622118 -2614 622354
rect -2378 622118 13198 622354
rect 13434 622118 13518 622354
rect 13754 622118 167826 622354
rect 168062 622118 168146 622354
rect 168382 622118 291590 622354
rect 291826 622118 291910 622354
rect 292146 622118 419826 622354
rect 420062 622118 420146 622354
rect 420382 622118 563826 622354
rect 564062 622118 564146 622354
rect 564382 622118 582326 622354
rect 582562 622118 582646 622354
rect 582882 622118 586302 622354
rect 586538 622118 586622 622354
rect 586858 622118 592650 622354
rect -8726 622034 592650 622118
rect -8726 621798 -2934 622034
rect -2698 621798 -2614 622034
rect -2378 621798 13198 622034
rect 13434 621798 13518 622034
rect 13754 621798 167826 622034
rect 168062 621798 168146 622034
rect 168382 621798 291590 622034
rect 291826 621798 291910 622034
rect 292146 621798 419826 622034
rect 420062 621798 420146 622034
rect 420382 621798 563826 622034
rect 564062 621798 564146 622034
rect 564382 621798 582326 622034
rect 582562 621798 582646 622034
rect 582882 621798 586302 622034
rect 586538 621798 586622 622034
rect 586858 621798 592650 622034
rect -8726 621766 592650 621798
rect -8726 617854 592650 617886
rect -8726 617618 -1974 617854
rect -1738 617618 -1654 617854
rect -1418 617618 5826 617854
rect 6062 617618 6146 617854
rect 6382 617618 173094 617854
rect 173330 617618 173414 617854
rect 173650 617618 293826 617854
rect 294062 617618 294146 617854
rect 294382 617618 401826 617854
rect 402062 617618 402146 617854
rect 402382 617618 570350 617854
rect 570586 617618 570670 617854
rect 570906 617618 585342 617854
rect 585578 617618 585662 617854
rect 585898 617618 592650 617854
rect -8726 617534 592650 617618
rect -8726 617298 -1974 617534
rect -1738 617298 -1654 617534
rect -1418 617298 5826 617534
rect 6062 617298 6146 617534
rect 6382 617298 173094 617534
rect 173330 617298 173414 617534
rect 173650 617298 293826 617534
rect 294062 617298 294146 617534
rect 294382 617298 401826 617534
rect 402062 617298 402146 617534
rect 402382 617298 570350 617534
rect 570586 617298 570670 617534
rect 570906 617298 585342 617534
rect 585578 617298 585662 617534
rect 585898 617298 592650 617534
rect -8726 617266 592650 617298
rect -8726 586354 592650 586386
rect -8726 586118 -2934 586354
rect -2698 586118 -2614 586354
rect -2378 586118 23826 586354
rect 24062 586118 24146 586354
rect 24382 586118 59826 586354
rect 60062 586118 60146 586354
rect 60382 586118 95826 586354
rect 96062 586118 96146 586354
rect 96382 586118 131826 586354
rect 132062 586118 132146 586354
rect 132382 586118 167826 586354
rect 168062 586118 168146 586354
rect 168382 586118 203826 586354
rect 204062 586118 204146 586354
rect 204382 586118 239826 586354
rect 240062 586118 240146 586354
rect 240382 586118 275826 586354
rect 276062 586118 276146 586354
rect 276382 586118 311826 586354
rect 312062 586118 312146 586354
rect 312382 586118 347826 586354
rect 348062 586118 348146 586354
rect 348382 586118 383826 586354
rect 384062 586118 384146 586354
rect 384382 586118 419826 586354
rect 420062 586118 420146 586354
rect 420382 586118 455826 586354
rect 456062 586118 456146 586354
rect 456382 586118 491826 586354
rect 492062 586118 492146 586354
rect 492382 586118 527826 586354
rect 528062 586118 528146 586354
rect 528382 586118 563826 586354
rect 564062 586118 564146 586354
rect 564382 586118 582326 586354
rect 582562 586118 582646 586354
rect 582882 586118 586302 586354
rect 586538 586118 586622 586354
rect 586858 586118 592650 586354
rect -8726 586034 592650 586118
rect -8726 585798 -2934 586034
rect -2698 585798 -2614 586034
rect -2378 585798 23826 586034
rect 24062 585798 24146 586034
rect 24382 585798 59826 586034
rect 60062 585798 60146 586034
rect 60382 585798 95826 586034
rect 96062 585798 96146 586034
rect 96382 585798 131826 586034
rect 132062 585798 132146 586034
rect 132382 585798 167826 586034
rect 168062 585798 168146 586034
rect 168382 585798 203826 586034
rect 204062 585798 204146 586034
rect 204382 585798 239826 586034
rect 240062 585798 240146 586034
rect 240382 585798 275826 586034
rect 276062 585798 276146 586034
rect 276382 585798 311826 586034
rect 312062 585798 312146 586034
rect 312382 585798 347826 586034
rect 348062 585798 348146 586034
rect 348382 585798 383826 586034
rect 384062 585798 384146 586034
rect 384382 585798 419826 586034
rect 420062 585798 420146 586034
rect 420382 585798 455826 586034
rect 456062 585798 456146 586034
rect 456382 585798 491826 586034
rect 492062 585798 492146 586034
rect 492382 585798 527826 586034
rect 528062 585798 528146 586034
rect 528382 585798 563826 586034
rect 564062 585798 564146 586034
rect 564382 585798 582326 586034
rect 582562 585798 582646 586034
rect 582882 585798 586302 586034
rect 586538 585798 586622 586034
rect 586858 585798 592650 586034
rect -8726 585766 592650 585798
rect -8726 581854 592650 581886
rect -8726 581618 -1974 581854
rect -1738 581618 -1654 581854
rect -1418 581618 5826 581854
rect 6062 581618 6146 581854
rect 6382 581618 41826 581854
rect 42062 581618 42146 581854
rect 42382 581618 77826 581854
rect 78062 581618 78146 581854
rect 78382 581618 113826 581854
rect 114062 581618 114146 581854
rect 114382 581618 149826 581854
rect 150062 581618 150146 581854
rect 150382 581618 185826 581854
rect 186062 581618 186146 581854
rect 186382 581618 221826 581854
rect 222062 581618 222146 581854
rect 222382 581618 257826 581854
rect 258062 581618 258146 581854
rect 258382 581618 293826 581854
rect 294062 581618 294146 581854
rect 294382 581618 329826 581854
rect 330062 581618 330146 581854
rect 330382 581618 365826 581854
rect 366062 581618 366146 581854
rect 366382 581618 401826 581854
rect 402062 581618 402146 581854
rect 402382 581618 437826 581854
rect 438062 581618 438146 581854
rect 438382 581618 473826 581854
rect 474062 581618 474146 581854
rect 474382 581618 509826 581854
rect 510062 581618 510146 581854
rect 510382 581618 545826 581854
rect 546062 581618 546146 581854
rect 546382 581618 585342 581854
rect 585578 581618 585662 581854
rect 585898 581618 592650 581854
rect -8726 581534 592650 581618
rect -8726 581298 -1974 581534
rect -1738 581298 -1654 581534
rect -1418 581298 5826 581534
rect 6062 581298 6146 581534
rect 6382 581298 41826 581534
rect 42062 581298 42146 581534
rect 42382 581298 77826 581534
rect 78062 581298 78146 581534
rect 78382 581298 113826 581534
rect 114062 581298 114146 581534
rect 114382 581298 149826 581534
rect 150062 581298 150146 581534
rect 150382 581298 185826 581534
rect 186062 581298 186146 581534
rect 186382 581298 221826 581534
rect 222062 581298 222146 581534
rect 222382 581298 257826 581534
rect 258062 581298 258146 581534
rect 258382 581298 293826 581534
rect 294062 581298 294146 581534
rect 294382 581298 329826 581534
rect 330062 581298 330146 581534
rect 330382 581298 365826 581534
rect 366062 581298 366146 581534
rect 366382 581298 401826 581534
rect 402062 581298 402146 581534
rect 402382 581298 437826 581534
rect 438062 581298 438146 581534
rect 438382 581298 473826 581534
rect 474062 581298 474146 581534
rect 474382 581298 509826 581534
rect 510062 581298 510146 581534
rect 510382 581298 545826 581534
rect 546062 581298 546146 581534
rect 546382 581298 585342 581534
rect 585578 581298 585662 581534
rect 585898 581298 592650 581534
rect -8726 581266 592650 581298
rect -8726 550354 592650 550386
rect -8726 550118 -2934 550354
rect -2698 550118 -2614 550354
rect -2378 550118 13198 550354
rect 13434 550118 13518 550354
rect 13754 550118 167826 550354
rect 168062 550118 168146 550354
rect 168382 550118 203826 550354
rect 204062 550118 204146 550354
rect 204382 550118 239826 550354
rect 240062 550118 240146 550354
rect 240382 550118 275826 550354
rect 276062 550118 276146 550354
rect 276382 550118 311826 550354
rect 312062 550118 312146 550354
rect 312382 550118 347826 550354
rect 348062 550118 348146 550354
rect 348382 550118 383826 550354
rect 384062 550118 384146 550354
rect 384382 550118 419826 550354
rect 420062 550118 420146 550354
rect 420382 550118 563826 550354
rect 564062 550118 564146 550354
rect 564382 550118 582326 550354
rect 582562 550118 582646 550354
rect 582882 550118 586302 550354
rect 586538 550118 586622 550354
rect 586858 550118 592650 550354
rect -8726 550034 592650 550118
rect -8726 549798 -2934 550034
rect -2698 549798 -2614 550034
rect -2378 549798 13198 550034
rect 13434 549798 13518 550034
rect 13754 549798 167826 550034
rect 168062 549798 168146 550034
rect 168382 549798 203826 550034
rect 204062 549798 204146 550034
rect 204382 549798 239826 550034
rect 240062 549798 240146 550034
rect 240382 549798 275826 550034
rect 276062 549798 276146 550034
rect 276382 549798 311826 550034
rect 312062 549798 312146 550034
rect 312382 549798 347826 550034
rect 348062 549798 348146 550034
rect 348382 549798 383826 550034
rect 384062 549798 384146 550034
rect 384382 549798 419826 550034
rect 420062 549798 420146 550034
rect 420382 549798 563826 550034
rect 564062 549798 564146 550034
rect 564382 549798 582326 550034
rect 582562 549798 582646 550034
rect 582882 549798 586302 550034
rect 586538 549798 586622 550034
rect 586858 549798 592650 550034
rect -8726 549766 592650 549798
rect -8726 545854 592650 545886
rect -8726 545618 -1974 545854
rect -1738 545618 -1654 545854
rect -1418 545618 5826 545854
rect 6062 545618 6146 545854
rect 6382 545618 185826 545854
rect 186062 545618 186146 545854
rect 186382 545618 221826 545854
rect 222062 545618 222146 545854
rect 222382 545618 257826 545854
rect 258062 545618 258146 545854
rect 258382 545618 293826 545854
rect 294062 545618 294146 545854
rect 294382 545618 329826 545854
rect 330062 545618 330146 545854
rect 330382 545618 365826 545854
rect 366062 545618 366146 545854
rect 366382 545618 401826 545854
rect 402062 545618 402146 545854
rect 402382 545618 570350 545854
rect 570586 545618 570670 545854
rect 570906 545618 585342 545854
rect 585578 545618 585662 545854
rect 585898 545618 592650 545854
rect -8726 545534 592650 545618
rect -8726 545298 -1974 545534
rect -1738 545298 -1654 545534
rect -1418 545298 5826 545534
rect 6062 545298 6146 545534
rect 6382 545298 185826 545534
rect 186062 545298 186146 545534
rect 186382 545298 221826 545534
rect 222062 545298 222146 545534
rect 222382 545298 257826 545534
rect 258062 545298 258146 545534
rect 258382 545298 293826 545534
rect 294062 545298 294146 545534
rect 294382 545298 329826 545534
rect 330062 545298 330146 545534
rect 330382 545298 365826 545534
rect 366062 545298 366146 545534
rect 366382 545298 401826 545534
rect 402062 545298 402146 545534
rect 402382 545298 570350 545534
rect 570586 545298 570670 545534
rect 570906 545298 585342 545534
rect 585578 545298 585662 545534
rect 585898 545298 592650 545534
rect -8726 545266 592650 545298
rect -8726 514354 592650 514386
rect -8726 514118 -2934 514354
rect -2698 514118 -2614 514354
rect -2378 514118 13198 514354
rect 13434 514118 13518 514354
rect 13754 514118 167826 514354
rect 168062 514118 168146 514354
rect 168382 514118 203826 514354
rect 204062 514118 204146 514354
rect 204382 514118 239826 514354
rect 240062 514118 240146 514354
rect 240382 514118 275826 514354
rect 276062 514118 276146 514354
rect 276382 514118 311826 514354
rect 312062 514118 312146 514354
rect 312382 514118 347826 514354
rect 348062 514118 348146 514354
rect 348382 514118 383826 514354
rect 384062 514118 384146 514354
rect 384382 514118 419826 514354
rect 420062 514118 420146 514354
rect 420382 514118 563826 514354
rect 564062 514118 564146 514354
rect 564382 514118 582326 514354
rect 582562 514118 582646 514354
rect 582882 514118 586302 514354
rect 586538 514118 586622 514354
rect 586858 514118 592650 514354
rect -8726 514034 592650 514118
rect -8726 513798 -2934 514034
rect -2698 513798 -2614 514034
rect -2378 513798 13198 514034
rect 13434 513798 13518 514034
rect 13754 513798 167826 514034
rect 168062 513798 168146 514034
rect 168382 513798 203826 514034
rect 204062 513798 204146 514034
rect 204382 513798 239826 514034
rect 240062 513798 240146 514034
rect 240382 513798 275826 514034
rect 276062 513798 276146 514034
rect 276382 513798 311826 514034
rect 312062 513798 312146 514034
rect 312382 513798 347826 514034
rect 348062 513798 348146 514034
rect 348382 513798 383826 514034
rect 384062 513798 384146 514034
rect 384382 513798 419826 514034
rect 420062 513798 420146 514034
rect 420382 513798 563826 514034
rect 564062 513798 564146 514034
rect 564382 513798 582326 514034
rect 582562 513798 582646 514034
rect 582882 513798 586302 514034
rect 586538 513798 586622 514034
rect 586858 513798 592650 514034
rect -8726 513766 592650 513798
rect -8726 509854 592650 509886
rect -8726 509618 -1974 509854
rect -1738 509618 -1654 509854
rect -1418 509618 5826 509854
rect 6062 509618 6146 509854
rect 6382 509618 185826 509854
rect 186062 509618 186146 509854
rect 186382 509618 221826 509854
rect 222062 509618 222146 509854
rect 222382 509618 257826 509854
rect 258062 509618 258146 509854
rect 258382 509618 293826 509854
rect 294062 509618 294146 509854
rect 294382 509618 329826 509854
rect 330062 509618 330146 509854
rect 330382 509618 365826 509854
rect 366062 509618 366146 509854
rect 366382 509618 401826 509854
rect 402062 509618 402146 509854
rect 402382 509618 570350 509854
rect 570586 509618 570670 509854
rect 570906 509618 585342 509854
rect 585578 509618 585662 509854
rect 585898 509618 592650 509854
rect -8726 509534 592650 509618
rect -8726 509298 -1974 509534
rect -1738 509298 -1654 509534
rect -1418 509298 5826 509534
rect 6062 509298 6146 509534
rect 6382 509298 185826 509534
rect 186062 509298 186146 509534
rect 186382 509298 221826 509534
rect 222062 509298 222146 509534
rect 222382 509298 257826 509534
rect 258062 509298 258146 509534
rect 258382 509298 293826 509534
rect 294062 509298 294146 509534
rect 294382 509298 329826 509534
rect 330062 509298 330146 509534
rect 330382 509298 365826 509534
rect 366062 509298 366146 509534
rect 366382 509298 401826 509534
rect 402062 509298 402146 509534
rect 402382 509298 570350 509534
rect 570586 509298 570670 509534
rect 570906 509298 585342 509534
rect 585578 509298 585662 509534
rect 585898 509298 592650 509534
rect -8726 509266 592650 509298
rect -8726 478354 592650 478386
rect -8726 478118 -2934 478354
rect -2698 478118 -2614 478354
rect -2378 478118 23826 478354
rect 24062 478118 24146 478354
rect 24382 478118 59826 478354
rect 60062 478118 60146 478354
rect 60382 478118 95826 478354
rect 96062 478118 96146 478354
rect 96382 478118 131826 478354
rect 132062 478118 132146 478354
rect 132382 478118 167826 478354
rect 168062 478118 168146 478354
rect 168382 478118 203826 478354
rect 204062 478118 204146 478354
rect 204382 478118 239826 478354
rect 240062 478118 240146 478354
rect 240382 478118 275826 478354
rect 276062 478118 276146 478354
rect 276382 478118 311826 478354
rect 312062 478118 312146 478354
rect 312382 478118 347826 478354
rect 348062 478118 348146 478354
rect 348382 478118 383826 478354
rect 384062 478118 384146 478354
rect 384382 478118 419826 478354
rect 420062 478118 420146 478354
rect 420382 478118 455826 478354
rect 456062 478118 456146 478354
rect 456382 478118 491826 478354
rect 492062 478118 492146 478354
rect 492382 478118 527826 478354
rect 528062 478118 528146 478354
rect 528382 478118 563826 478354
rect 564062 478118 564146 478354
rect 564382 478118 582326 478354
rect 582562 478118 582646 478354
rect 582882 478118 586302 478354
rect 586538 478118 586622 478354
rect 586858 478118 592650 478354
rect -8726 478034 592650 478118
rect -8726 477798 -2934 478034
rect -2698 477798 -2614 478034
rect -2378 477798 23826 478034
rect 24062 477798 24146 478034
rect 24382 477798 59826 478034
rect 60062 477798 60146 478034
rect 60382 477798 95826 478034
rect 96062 477798 96146 478034
rect 96382 477798 131826 478034
rect 132062 477798 132146 478034
rect 132382 477798 167826 478034
rect 168062 477798 168146 478034
rect 168382 477798 203826 478034
rect 204062 477798 204146 478034
rect 204382 477798 239826 478034
rect 240062 477798 240146 478034
rect 240382 477798 275826 478034
rect 276062 477798 276146 478034
rect 276382 477798 311826 478034
rect 312062 477798 312146 478034
rect 312382 477798 347826 478034
rect 348062 477798 348146 478034
rect 348382 477798 383826 478034
rect 384062 477798 384146 478034
rect 384382 477798 419826 478034
rect 420062 477798 420146 478034
rect 420382 477798 455826 478034
rect 456062 477798 456146 478034
rect 456382 477798 491826 478034
rect 492062 477798 492146 478034
rect 492382 477798 527826 478034
rect 528062 477798 528146 478034
rect 528382 477798 563826 478034
rect 564062 477798 564146 478034
rect 564382 477798 582326 478034
rect 582562 477798 582646 478034
rect 582882 477798 586302 478034
rect 586538 477798 586622 478034
rect 586858 477798 592650 478034
rect -8726 477766 592650 477798
rect -8726 473854 592650 473886
rect -8726 473618 -1974 473854
rect -1738 473618 -1654 473854
rect -1418 473618 5826 473854
rect 6062 473618 6146 473854
rect 6382 473618 41826 473854
rect 42062 473618 42146 473854
rect 42382 473618 77826 473854
rect 78062 473618 78146 473854
rect 78382 473618 113826 473854
rect 114062 473618 114146 473854
rect 114382 473618 149826 473854
rect 150062 473618 150146 473854
rect 150382 473618 185826 473854
rect 186062 473618 186146 473854
rect 186382 473618 221826 473854
rect 222062 473618 222146 473854
rect 222382 473618 257826 473854
rect 258062 473618 258146 473854
rect 258382 473618 293826 473854
rect 294062 473618 294146 473854
rect 294382 473618 329826 473854
rect 330062 473618 330146 473854
rect 330382 473618 365826 473854
rect 366062 473618 366146 473854
rect 366382 473618 401826 473854
rect 402062 473618 402146 473854
rect 402382 473618 437826 473854
rect 438062 473618 438146 473854
rect 438382 473618 473826 473854
rect 474062 473618 474146 473854
rect 474382 473618 509826 473854
rect 510062 473618 510146 473854
rect 510382 473618 545826 473854
rect 546062 473618 546146 473854
rect 546382 473618 585342 473854
rect 585578 473618 585662 473854
rect 585898 473618 592650 473854
rect -8726 473534 592650 473618
rect -8726 473298 -1974 473534
rect -1738 473298 -1654 473534
rect -1418 473298 5826 473534
rect 6062 473298 6146 473534
rect 6382 473298 41826 473534
rect 42062 473298 42146 473534
rect 42382 473298 77826 473534
rect 78062 473298 78146 473534
rect 78382 473298 113826 473534
rect 114062 473298 114146 473534
rect 114382 473298 149826 473534
rect 150062 473298 150146 473534
rect 150382 473298 185826 473534
rect 186062 473298 186146 473534
rect 186382 473298 221826 473534
rect 222062 473298 222146 473534
rect 222382 473298 257826 473534
rect 258062 473298 258146 473534
rect 258382 473298 293826 473534
rect 294062 473298 294146 473534
rect 294382 473298 329826 473534
rect 330062 473298 330146 473534
rect 330382 473298 365826 473534
rect 366062 473298 366146 473534
rect 366382 473298 401826 473534
rect 402062 473298 402146 473534
rect 402382 473298 437826 473534
rect 438062 473298 438146 473534
rect 438382 473298 473826 473534
rect 474062 473298 474146 473534
rect 474382 473298 509826 473534
rect 510062 473298 510146 473534
rect 510382 473298 545826 473534
rect 546062 473298 546146 473534
rect 546382 473298 585342 473534
rect 585578 473298 585662 473534
rect 585898 473298 592650 473534
rect -8726 473266 592650 473298
rect -8726 442354 592650 442386
rect -8726 442118 -2934 442354
rect -2698 442118 -2614 442354
rect -2378 442118 13198 442354
rect 13434 442118 13518 442354
rect 13754 442118 167826 442354
rect 168062 442118 168146 442354
rect 168382 442118 203826 442354
rect 204062 442118 204146 442354
rect 204382 442118 239826 442354
rect 240062 442118 240146 442354
rect 240382 442118 275826 442354
rect 276062 442118 276146 442354
rect 276382 442118 311826 442354
rect 312062 442118 312146 442354
rect 312382 442118 347826 442354
rect 348062 442118 348146 442354
rect 348382 442118 383826 442354
rect 384062 442118 384146 442354
rect 384382 442118 419826 442354
rect 420062 442118 420146 442354
rect 420382 442118 563826 442354
rect 564062 442118 564146 442354
rect 564382 442118 582326 442354
rect 582562 442118 582646 442354
rect 582882 442118 586302 442354
rect 586538 442118 586622 442354
rect 586858 442118 592650 442354
rect -8726 442034 592650 442118
rect -8726 441798 -2934 442034
rect -2698 441798 -2614 442034
rect -2378 441798 13198 442034
rect 13434 441798 13518 442034
rect 13754 441798 167826 442034
rect 168062 441798 168146 442034
rect 168382 441798 203826 442034
rect 204062 441798 204146 442034
rect 204382 441798 239826 442034
rect 240062 441798 240146 442034
rect 240382 441798 275826 442034
rect 276062 441798 276146 442034
rect 276382 441798 311826 442034
rect 312062 441798 312146 442034
rect 312382 441798 347826 442034
rect 348062 441798 348146 442034
rect 348382 441798 383826 442034
rect 384062 441798 384146 442034
rect 384382 441798 419826 442034
rect 420062 441798 420146 442034
rect 420382 441798 563826 442034
rect 564062 441798 564146 442034
rect 564382 441798 582326 442034
rect 582562 441798 582646 442034
rect 582882 441798 586302 442034
rect 586538 441798 586622 442034
rect 586858 441798 592650 442034
rect -8726 441766 592650 441798
rect -8726 437854 592650 437886
rect -8726 437618 -1974 437854
rect -1738 437618 -1654 437854
rect -1418 437618 5826 437854
rect 6062 437618 6146 437854
rect 6382 437618 185826 437854
rect 186062 437618 186146 437854
rect 186382 437618 221826 437854
rect 222062 437618 222146 437854
rect 222382 437618 257826 437854
rect 258062 437618 258146 437854
rect 258382 437618 293826 437854
rect 294062 437618 294146 437854
rect 294382 437618 329826 437854
rect 330062 437618 330146 437854
rect 330382 437618 365826 437854
rect 366062 437618 366146 437854
rect 366382 437618 401826 437854
rect 402062 437618 402146 437854
rect 402382 437618 570350 437854
rect 570586 437618 570670 437854
rect 570906 437618 585342 437854
rect 585578 437618 585662 437854
rect 585898 437618 592650 437854
rect -8726 437534 592650 437618
rect -8726 437298 -1974 437534
rect -1738 437298 -1654 437534
rect -1418 437298 5826 437534
rect 6062 437298 6146 437534
rect 6382 437298 185826 437534
rect 186062 437298 186146 437534
rect 186382 437298 221826 437534
rect 222062 437298 222146 437534
rect 222382 437298 257826 437534
rect 258062 437298 258146 437534
rect 258382 437298 293826 437534
rect 294062 437298 294146 437534
rect 294382 437298 329826 437534
rect 330062 437298 330146 437534
rect 330382 437298 365826 437534
rect 366062 437298 366146 437534
rect 366382 437298 401826 437534
rect 402062 437298 402146 437534
rect 402382 437298 570350 437534
rect 570586 437298 570670 437534
rect 570906 437298 585342 437534
rect 585578 437298 585662 437534
rect 585898 437298 592650 437534
rect -8726 437266 592650 437298
rect -8726 406354 592650 406386
rect -8726 406118 -2934 406354
rect -2698 406118 -2614 406354
rect -2378 406118 13198 406354
rect 13434 406118 13518 406354
rect 13754 406118 167826 406354
rect 168062 406118 168146 406354
rect 168382 406118 203826 406354
rect 204062 406118 204146 406354
rect 204382 406118 239826 406354
rect 240062 406118 240146 406354
rect 240382 406118 275826 406354
rect 276062 406118 276146 406354
rect 276382 406118 311826 406354
rect 312062 406118 312146 406354
rect 312382 406118 347826 406354
rect 348062 406118 348146 406354
rect 348382 406118 383826 406354
rect 384062 406118 384146 406354
rect 384382 406118 419826 406354
rect 420062 406118 420146 406354
rect 420382 406118 563826 406354
rect 564062 406118 564146 406354
rect 564382 406118 582326 406354
rect 582562 406118 582646 406354
rect 582882 406118 586302 406354
rect 586538 406118 586622 406354
rect 586858 406118 592650 406354
rect -8726 406034 592650 406118
rect -8726 405798 -2934 406034
rect -2698 405798 -2614 406034
rect -2378 405798 13198 406034
rect 13434 405798 13518 406034
rect 13754 405798 167826 406034
rect 168062 405798 168146 406034
rect 168382 405798 203826 406034
rect 204062 405798 204146 406034
rect 204382 405798 239826 406034
rect 240062 405798 240146 406034
rect 240382 405798 275826 406034
rect 276062 405798 276146 406034
rect 276382 405798 311826 406034
rect 312062 405798 312146 406034
rect 312382 405798 347826 406034
rect 348062 405798 348146 406034
rect 348382 405798 383826 406034
rect 384062 405798 384146 406034
rect 384382 405798 419826 406034
rect 420062 405798 420146 406034
rect 420382 405798 563826 406034
rect 564062 405798 564146 406034
rect 564382 405798 582326 406034
rect 582562 405798 582646 406034
rect 582882 405798 586302 406034
rect 586538 405798 586622 406034
rect 586858 405798 592650 406034
rect -8726 405766 592650 405798
rect -8726 401854 592650 401886
rect -8726 401618 -1974 401854
rect -1738 401618 -1654 401854
rect -1418 401618 5826 401854
rect 6062 401618 6146 401854
rect 6382 401618 185826 401854
rect 186062 401618 186146 401854
rect 186382 401618 221826 401854
rect 222062 401618 222146 401854
rect 222382 401618 257826 401854
rect 258062 401618 258146 401854
rect 258382 401618 293826 401854
rect 294062 401618 294146 401854
rect 294382 401618 329826 401854
rect 330062 401618 330146 401854
rect 330382 401618 365826 401854
rect 366062 401618 366146 401854
rect 366382 401618 401826 401854
rect 402062 401618 402146 401854
rect 402382 401618 570350 401854
rect 570586 401618 570670 401854
rect 570906 401618 585342 401854
rect 585578 401618 585662 401854
rect 585898 401618 592650 401854
rect -8726 401534 592650 401618
rect -8726 401298 -1974 401534
rect -1738 401298 -1654 401534
rect -1418 401298 5826 401534
rect 6062 401298 6146 401534
rect 6382 401298 185826 401534
rect 186062 401298 186146 401534
rect 186382 401298 221826 401534
rect 222062 401298 222146 401534
rect 222382 401298 257826 401534
rect 258062 401298 258146 401534
rect 258382 401298 293826 401534
rect 294062 401298 294146 401534
rect 294382 401298 329826 401534
rect 330062 401298 330146 401534
rect 330382 401298 365826 401534
rect 366062 401298 366146 401534
rect 366382 401298 401826 401534
rect 402062 401298 402146 401534
rect 402382 401298 570350 401534
rect 570586 401298 570670 401534
rect 570906 401298 585342 401534
rect 585578 401298 585662 401534
rect 585898 401298 592650 401534
rect -8726 401266 592650 401298
rect -8726 370354 592650 370386
rect -8726 370118 -2934 370354
rect -2698 370118 -2614 370354
rect -2378 370118 13198 370354
rect 13434 370118 13518 370354
rect 13754 370118 167826 370354
rect 168062 370118 168146 370354
rect 168382 370118 203826 370354
rect 204062 370118 204146 370354
rect 204382 370118 239826 370354
rect 240062 370118 240146 370354
rect 240382 370118 275826 370354
rect 276062 370118 276146 370354
rect 276382 370118 311826 370354
rect 312062 370118 312146 370354
rect 312382 370118 347826 370354
rect 348062 370118 348146 370354
rect 348382 370118 383826 370354
rect 384062 370118 384146 370354
rect 384382 370118 419826 370354
rect 420062 370118 420146 370354
rect 420382 370118 563826 370354
rect 564062 370118 564146 370354
rect 564382 370118 582326 370354
rect 582562 370118 582646 370354
rect 582882 370118 586302 370354
rect 586538 370118 586622 370354
rect 586858 370118 592650 370354
rect -8726 370034 592650 370118
rect -8726 369798 -2934 370034
rect -2698 369798 -2614 370034
rect -2378 369798 13198 370034
rect 13434 369798 13518 370034
rect 13754 369798 167826 370034
rect 168062 369798 168146 370034
rect 168382 369798 203826 370034
rect 204062 369798 204146 370034
rect 204382 369798 239826 370034
rect 240062 369798 240146 370034
rect 240382 369798 275826 370034
rect 276062 369798 276146 370034
rect 276382 369798 311826 370034
rect 312062 369798 312146 370034
rect 312382 369798 347826 370034
rect 348062 369798 348146 370034
rect 348382 369798 383826 370034
rect 384062 369798 384146 370034
rect 384382 369798 419826 370034
rect 420062 369798 420146 370034
rect 420382 369798 563826 370034
rect 564062 369798 564146 370034
rect 564382 369798 582326 370034
rect 582562 369798 582646 370034
rect 582882 369798 586302 370034
rect 586538 369798 586622 370034
rect 586858 369798 592650 370034
rect -8726 369766 592650 369798
rect -8726 365854 592650 365886
rect -8726 365618 -1974 365854
rect -1738 365618 -1654 365854
rect -1418 365618 5826 365854
rect 6062 365618 6146 365854
rect 6382 365618 41826 365854
rect 42062 365618 42146 365854
rect 42382 365618 77826 365854
rect 78062 365618 78146 365854
rect 78382 365618 113826 365854
rect 114062 365618 114146 365854
rect 114382 365618 149826 365854
rect 150062 365618 150146 365854
rect 150382 365618 185826 365854
rect 186062 365618 186146 365854
rect 186382 365618 221826 365854
rect 222062 365618 222146 365854
rect 222382 365618 257826 365854
rect 258062 365618 258146 365854
rect 258382 365618 293826 365854
rect 294062 365618 294146 365854
rect 294382 365618 329826 365854
rect 330062 365618 330146 365854
rect 330382 365618 365826 365854
rect 366062 365618 366146 365854
rect 366382 365618 401826 365854
rect 402062 365618 402146 365854
rect 402382 365618 437826 365854
rect 438062 365618 438146 365854
rect 438382 365618 473826 365854
rect 474062 365618 474146 365854
rect 474382 365618 509826 365854
rect 510062 365618 510146 365854
rect 510382 365618 545826 365854
rect 546062 365618 546146 365854
rect 546382 365618 585342 365854
rect 585578 365618 585662 365854
rect 585898 365618 592650 365854
rect -8726 365534 592650 365618
rect -8726 365298 -1974 365534
rect -1738 365298 -1654 365534
rect -1418 365298 5826 365534
rect 6062 365298 6146 365534
rect 6382 365298 41826 365534
rect 42062 365298 42146 365534
rect 42382 365298 77826 365534
rect 78062 365298 78146 365534
rect 78382 365298 113826 365534
rect 114062 365298 114146 365534
rect 114382 365298 149826 365534
rect 150062 365298 150146 365534
rect 150382 365298 185826 365534
rect 186062 365298 186146 365534
rect 186382 365298 221826 365534
rect 222062 365298 222146 365534
rect 222382 365298 257826 365534
rect 258062 365298 258146 365534
rect 258382 365298 293826 365534
rect 294062 365298 294146 365534
rect 294382 365298 329826 365534
rect 330062 365298 330146 365534
rect 330382 365298 365826 365534
rect 366062 365298 366146 365534
rect 366382 365298 401826 365534
rect 402062 365298 402146 365534
rect 402382 365298 437826 365534
rect 438062 365298 438146 365534
rect 438382 365298 473826 365534
rect 474062 365298 474146 365534
rect 474382 365298 509826 365534
rect 510062 365298 510146 365534
rect 510382 365298 545826 365534
rect 546062 365298 546146 365534
rect 546382 365298 585342 365534
rect 585578 365298 585662 365534
rect 585898 365298 592650 365534
rect -8726 365266 592650 365298
rect -8726 334354 592650 334386
rect -8726 334118 -2934 334354
rect -2698 334118 -2614 334354
rect -2378 334118 13198 334354
rect 13434 334118 13518 334354
rect 13754 334118 167826 334354
rect 168062 334118 168146 334354
rect 168382 334118 203826 334354
rect 204062 334118 204146 334354
rect 204382 334118 239826 334354
rect 240062 334118 240146 334354
rect 240382 334118 275826 334354
rect 276062 334118 276146 334354
rect 276382 334118 311826 334354
rect 312062 334118 312146 334354
rect 312382 334118 347826 334354
rect 348062 334118 348146 334354
rect 348382 334118 383826 334354
rect 384062 334118 384146 334354
rect 384382 334118 419826 334354
rect 420062 334118 420146 334354
rect 420382 334118 563826 334354
rect 564062 334118 564146 334354
rect 564382 334118 582326 334354
rect 582562 334118 582646 334354
rect 582882 334118 586302 334354
rect 586538 334118 586622 334354
rect 586858 334118 592650 334354
rect -8726 334034 592650 334118
rect -8726 333798 -2934 334034
rect -2698 333798 -2614 334034
rect -2378 333798 13198 334034
rect 13434 333798 13518 334034
rect 13754 333798 167826 334034
rect 168062 333798 168146 334034
rect 168382 333798 203826 334034
rect 204062 333798 204146 334034
rect 204382 333798 239826 334034
rect 240062 333798 240146 334034
rect 240382 333798 275826 334034
rect 276062 333798 276146 334034
rect 276382 333798 311826 334034
rect 312062 333798 312146 334034
rect 312382 333798 347826 334034
rect 348062 333798 348146 334034
rect 348382 333798 383826 334034
rect 384062 333798 384146 334034
rect 384382 333798 419826 334034
rect 420062 333798 420146 334034
rect 420382 333798 563826 334034
rect 564062 333798 564146 334034
rect 564382 333798 582326 334034
rect 582562 333798 582646 334034
rect 582882 333798 586302 334034
rect 586538 333798 586622 334034
rect 586858 333798 592650 334034
rect -8726 333766 592650 333798
rect -8726 329854 592650 329886
rect -8726 329618 -1974 329854
rect -1738 329618 -1654 329854
rect -1418 329618 5826 329854
rect 6062 329618 6146 329854
rect 6382 329618 185826 329854
rect 186062 329618 186146 329854
rect 186382 329618 221826 329854
rect 222062 329618 222146 329854
rect 222382 329618 257826 329854
rect 258062 329618 258146 329854
rect 258382 329618 293826 329854
rect 294062 329618 294146 329854
rect 294382 329618 329826 329854
rect 330062 329618 330146 329854
rect 330382 329618 365826 329854
rect 366062 329618 366146 329854
rect 366382 329618 401826 329854
rect 402062 329618 402146 329854
rect 402382 329618 570350 329854
rect 570586 329618 570670 329854
rect 570906 329618 585342 329854
rect 585578 329618 585662 329854
rect 585898 329618 592650 329854
rect -8726 329534 592650 329618
rect -8726 329298 -1974 329534
rect -1738 329298 -1654 329534
rect -1418 329298 5826 329534
rect 6062 329298 6146 329534
rect 6382 329298 185826 329534
rect 186062 329298 186146 329534
rect 186382 329298 221826 329534
rect 222062 329298 222146 329534
rect 222382 329298 257826 329534
rect 258062 329298 258146 329534
rect 258382 329298 293826 329534
rect 294062 329298 294146 329534
rect 294382 329298 329826 329534
rect 330062 329298 330146 329534
rect 330382 329298 365826 329534
rect 366062 329298 366146 329534
rect 366382 329298 401826 329534
rect 402062 329298 402146 329534
rect 402382 329298 570350 329534
rect 570586 329298 570670 329534
rect 570906 329298 585342 329534
rect 585578 329298 585662 329534
rect 585898 329298 592650 329534
rect -8726 329266 592650 329298
rect -8726 298354 592650 298386
rect -8726 298118 -2934 298354
rect -2698 298118 -2614 298354
rect -2378 298118 13198 298354
rect 13434 298118 13518 298354
rect 13754 298118 167826 298354
rect 168062 298118 168146 298354
rect 168382 298118 203826 298354
rect 204062 298118 204146 298354
rect 204382 298118 239826 298354
rect 240062 298118 240146 298354
rect 240382 298118 275826 298354
rect 276062 298118 276146 298354
rect 276382 298118 311826 298354
rect 312062 298118 312146 298354
rect 312382 298118 347826 298354
rect 348062 298118 348146 298354
rect 348382 298118 383826 298354
rect 384062 298118 384146 298354
rect 384382 298118 419826 298354
rect 420062 298118 420146 298354
rect 420382 298118 563826 298354
rect 564062 298118 564146 298354
rect 564382 298118 582326 298354
rect 582562 298118 582646 298354
rect 582882 298118 586302 298354
rect 586538 298118 586622 298354
rect 586858 298118 592650 298354
rect -8726 298034 592650 298118
rect -8726 297798 -2934 298034
rect -2698 297798 -2614 298034
rect -2378 297798 13198 298034
rect 13434 297798 13518 298034
rect 13754 297798 167826 298034
rect 168062 297798 168146 298034
rect 168382 297798 203826 298034
rect 204062 297798 204146 298034
rect 204382 297798 239826 298034
rect 240062 297798 240146 298034
rect 240382 297798 275826 298034
rect 276062 297798 276146 298034
rect 276382 297798 311826 298034
rect 312062 297798 312146 298034
rect 312382 297798 347826 298034
rect 348062 297798 348146 298034
rect 348382 297798 383826 298034
rect 384062 297798 384146 298034
rect 384382 297798 419826 298034
rect 420062 297798 420146 298034
rect 420382 297798 563826 298034
rect 564062 297798 564146 298034
rect 564382 297798 582326 298034
rect 582562 297798 582646 298034
rect 582882 297798 586302 298034
rect 586538 297798 586622 298034
rect 586858 297798 592650 298034
rect -8726 297766 592650 297798
rect -8726 293854 592650 293886
rect -8726 293618 -1974 293854
rect -1738 293618 -1654 293854
rect -1418 293618 5826 293854
rect 6062 293618 6146 293854
rect 6382 293618 185826 293854
rect 186062 293618 186146 293854
rect 186382 293618 221826 293854
rect 222062 293618 222146 293854
rect 222382 293618 257826 293854
rect 258062 293618 258146 293854
rect 258382 293618 293826 293854
rect 294062 293618 294146 293854
rect 294382 293618 329826 293854
rect 330062 293618 330146 293854
rect 330382 293618 365826 293854
rect 366062 293618 366146 293854
rect 366382 293618 401826 293854
rect 402062 293618 402146 293854
rect 402382 293618 570350 293854
rect 570586 293618 570670 293854
rect 570906 293618 585342 293854
rect 585578 293618 585662 293854
rect 585898 293618 592650 293854
rect -8726 293534 592650 293618
rect -8726 293298 -1974 293534
rect -1738 293298 -1654 293534
rect -1418 293298 5826 293534
rect 6062 293298 6146 293534
rect 6382 293298 185826 293534
rect 186062 293298 186146 293534
rect 186382 293298 221826 293534
rect 222062 293298 222146 293534
rect 222382 293298 257826 293534
rect 258062 293298 258146 293534
rect 258382 293298 293826 293534
rect 294062 293298 294146 293534
rect 294382 293298 329826 293534
rect 330062 293298 330146 293534
rect 330382 293298 365826 293534
rect 366062 293298 366146 293534
rect 366382 293298 401826 293534
rect 402062 293298 402146 293534
rect 402382 293298 570350 293534
rect 570586 293298 570670 293534
rect 570906 293298 585342 293534
rect 585578 293298 585662 293534
rect 585898 293298 592650 293534
rect -8726 293266 592650 293298
rect -8726 262354 592650 262386
rect -8726 262118 -2934 262354
rect -2698 262118 -2614 262354
rect -2378 262118 13198 262354
rect 13434 262118 13518 262354
rect 13754 262118 167826 262354
rect 168062 262118 168146 262354
rect 168382 262118 203826 262354
rect 204062 262118 204146 262354
rect 204382 262118 239826 262354
rect 240062 262118 240146 262354
rect 240382 262118 275826 262354
rect 276062 262118 276146 262354
rect 276382 262118 311826 262354
rect 312062 262118 312146 262354
rect 312382 262118 347826 262354
rect 348062 262118 348146 262354
rect 348382 262118 383826 262354
rect 384062 262118 384146 262354
rect 384382 262118 419826 262354
rect 420062 262118 420146 262354
rect 420382 262118 563826 262354
rect 564062 262118 564146 262354
rect 564382 262118 582326 262354
rect 582562 262118 582646 262354
rect 582882 262118 586302 262354
rect 586538 262118 586622 262354
rect 586858 262118 592650 262354
rect -8726 262034 592650 262118
rect -8726 261798 -2934 262034
rect -2698 261798 -2614 262034
rect -2378 261798 13198 262034
rect 13434 261798 13518 262034
rect 13754 261798 167826 262034
rect 168062 261798 168146 262034
rect 168382 261798 203826 262034
rect 204062 261798 204146 262034
rect 204382 261798 239826 262034
rect 240062 261798 240146 262034
rect 240382 261798 275826 262034
rect 276062 261798 276146 262034
rect 276382 261798 311826 262034
rect 312062 261798 312146 262034
rect 312382 261798 347826 262034
rect 348062 261798 348146 262034
rect 348382 261798 383826 262034
rect 384062 261798 384146 262034
rect 384382 261798 419826 262034
rect 420062 261798 420146 262034
rect 420382 261798 563826 262034
rect 564062 261798 564146 262034
rect 564382 261798 582326 262034
rect 582562 261798 582646 262034
rect 582882 261798 586302 262034
rect 586538 261798 586622 262034
rect 586858 261798 592650 262034
rect -8726 261766 592650 261798
rect -8726 257854 592650 257886
rect -8726 257618 -1974 257854
rect -1738 257618 -1654 257854
rect -1418 257618 5826 257854
rect 6062 257618 6146 257854
rect 6382 257618 185826 257854
rect 186062 257618 186146 257854
rect 186382 257618 221826 257854
rect 222062 257618 222146 257854
rect 222382 257618 257826 257854
rect 258062 257618 258146 257854
rect 258382 257618 293826 257854
rect 294062 257618 294146 257854
rect 294382 257618 329826 257854
rect 330062 257618 330146 257854
rect 330382 257618 365826 257854
rect 366062 257618 366146 257854
rect 366382 257618 401826 257854
rect 402062 257618 402146 257854
rect 402382 257618 570350 257854
rect 570586 257618 570670 257854
rect 570906 257618 585342 257854
rect 585578 257618 585662 257854
rect 585898 257618 592650 257854
rect -8726 257534 592650 257618
rect -8726 257298 -1974 257534
rect -1738 257298 -1654 257534
rect -1418 257298 5826 257534
rect 6062 257298 6146 257534
rect 6382 257298 185826 257534
rect 186062 257298 186146 257534
rect 186382 257298 221826 257534
rect 222062 257298 222146 257534
rect 222382 257298 257826 257534
rect 258062 257298 258146 257534
rect 258382 257298 293826 257534
rect 294062 257298 294146 257534
rect 294382 257298 329826 257534
rect 330062 257298 330146 257534
rect 330382 257298 365826 257534
rect 366062 257298 366146 257534
rect 366382 257298 401826 257534
rect 402062 257298 402146 257534
rect 402382 257298 570350 257534
rect 570586 257298 570670 257534
rect 570906 257298 585342 257534
rect 585578 257298 585662 257534
rect 585898 257298 592650 257534
rect -8726 257266 592650 257298
rect -8726 226354 592650 226386
rect -8726 226118 -2934 226354
rect -2698 226118 -2614 226354
rect -2378 226118 23826 226354
rect 24062 226118 24146 226354
rect 24382 226118 59826 226354
rect 60062 226118 60146 226354
rect 60382 226118 95826 226354
rect 96062 226118 96146 226354
rect 96382 226118 131826 226354
rect 132062 226118 132146 226354
rect 132382 226118 167826 226354
rect 168062 226118 168146 226354
rect 168382 226118 203826 226354
rect 204062 226118 204146 226354
rect 204382 226118 239826 226354
rect 240062 226118 240146 226354
rect 240382 226118 275826 226354
rect 276062 226118 276146 226354
rect 276382 226118 311826 226354
rect 312062 226118 312146 226354
rect 312382 226118 347826 226354
rect 348062 226118 348146 226354
rect 348382 226118 383826 226354
rect 384062 226118 384146 226354
rect 384382 226118 419826 226354
rect 420062 226118 420146 226354
rect 420382 226118 455826 226354
rect 456062 226118 456146 226354
rect 456382 226118 491826 226354
rect 492062 226118 492146 226354
rect 492382 226118 527826 226354
rect 528062 226118 528146 226354
rect 528382 226118 563826 226354
rect 564062 226118 564146 226354
rect 564382 226118 582326 226354
rect 582562 226118 582646 226354
rect 582882 226118 586302 226354
rect 586538 226118 586622 226354
rect 586858 226118 592650 226354
rect -8726 226034 592650 226118
rect -8726 225798 -2934 226034
rect -2698 225798 -2614 226034
rect -2378 225798 23826 226034
rect 24062 225798 24146 226034
rect 24382 225798 59826 226034
rect 60062 225798 60146 226034
rect 60382 225798 95826 226034
rect 96062 225798 96146 226034
rect 96382 225798 131826 226034
rect 132062 225798 132146 226034
rect 132382 225798 167826 226034
rect 168062 225798 168146 226034
rect 168382 225798 203826 226034
rect 204062 225798 204146 226034
rect 204382 225798 239826 226034
rect 240062 225798 240146 226034
rect 240382 225798 275826 226034
rect 276062 225798 276146 226034
rect 276382 225798 311826 226034
rect 312062 225798 312146 226034
rect 312382 225798 347826 226034
rect 348062 225798 348146 226034
rect 348382 225798 383826 226034
rect 384062 225798 384146 226034
rect 384382 225798 419826 226034
rect 420062 225798 420146 226034
rect 420382 225798 455826 226034
rect 456062 225798 456146 226034
rect 456382 225798 491826 226034
rect 492062 225798 492146 226034
rect 492382 225798 527826 226034
rect 528062 225798 528146 226034
rect 528382 225798 563826 226034
rect 564062 225798 564146 226034
rect 564382 225798 582326 226034
rect 582562 225798 582646 226034
rect 582882 225798 586302 226034
rect 586538 225798 586622 226034
rect 586858 225798 592650 226034
rect -8726 225766 592650 225798
rect -8726 221854 592650 221886
rect -8726 221618 -1974 221854
rect -1738 221618 -1654 221854
rect -1418 221618 5826 221854
rect 6062 221618 6146 221854
rect 6382 221618 185826 221854
rect 186062 221618 186146 221854
rect 186382 221618 221826 221854
rect 222062 221618 222146 221854
rect 222382 221618 257826 221854
rect 258062 221618 258146 221854
rect 258382 221618 293826 221854
rect 294062 221618 294146 221854
rect 294382 221618 329826 221854
rect 330062 221618 330146 221854
rect 330382 221618 365826 221854
rect 366062 221618 366146 221854
rect 366382 221618 401826 221854
rect 402062 221618 402146 221854
rect 402382 221618 570350 221854
rect 570586 221618 570670 221854
rect 570906 221618 585342 221854
rect 585578 221618 585662 221854
rect 585898 221618 592650 221854
rect -8726 221534 592650 221618
rect -8726 221298 -1974 221534
rect -1738 221298 -1654 221534
rect -1418 221298 5826 221534
rect 6062 221298 6146 221534
rect 6382 221298 185826 221534
rect 186062 221298 186146 221534
rect 186382 221298 221826 221534
rect 222062 221298 222146 221534
rect 222382 221298 257826 221534
rect 258062 221298 258146 221534
rect 258382 221298 293826 221534
rect 294062 221298 294146 221534
rect 294382 221298 329826 221534
rect 330062 221298 330146 221534
rect 330382 221298 365826 221534
rect 366062 221298 366146 221534
rect 366382 221298 401826 221534
rect 402062 221298 402146 221534
rect 402382 221298 570350 221534
rect 570586 221298 570670 221534
rect 570906 221298 585342 221534
rect 585578 221298 585662 221534
rect 585898 221298 592650 221534
rect -8726 221266 592650 221298
rect -8726 190354 592650 190386
rect -8726 190118 -2934 190354
rect -2698 190118 -2614 190354
rect -2378 190118 13198 190354
rect 13434 190118 13518 190354
rect 13754 190118 167826 190354
rect 168062 190118 168146 190354
rect 168382 190118 203826 190354
rect 204062 190118 204146 190354
rect 204382 190118 239826 190354
rect 240062 190118 240146 190354
rect 240382 190118 275826 190354
rect 276062 190118 276146 190354
rect 276382 190118 311826 190354
rect 312062 190118 312146 190354
rect 312382 190118 347826 190354
rect 348062 190118 348146 190354
rect 348382 190118 383826 190354
rect 384062 190118 384146 190354
rect 384382 190118 419826 190354
rect 420062 190118 420146 190354
rect 420382 190118 563826 190354
rect 564062 190118 564146 190354
rect 564382 190118 582326 190354
rect 582562 190118 582646 190354
rect 582882 190118 586302 190354
rect 586538 190118 586622 190354
rect 586858 190118 592650 190354
rect -8726 190034 592650 190118
rect -8726 189798 -2934 190034
rect -2698 189798 -2614 190034
rect -2378 189798 13198 190034
rect 13434 189798 13518 190034
rect 13754 189798 167826 190034
rect 168062 189798 168146 190034
rect 168382 189798 203826 190034
rect 204062 189798 204146 190034
rect 204382 189798 239826 190034
rect 240062 189798 240146 190034
rect 240382 189798 275826 190034
rect 276062 189798 276146 190034
rect 276382 189798 311826 190034
rect 312062 189798 312146 190034
rect 312382 189798 347826 190034
rect 348062 189798 348146 190034
rect 348382 189798 383826 190034
rect 384062 189798 384146 190034
rect 384382 189798 419826 190034
rect 420062 189798 420146 190034
rect 420382 189798 563826 190034
rect 564062 189798 564146 190034
rect 564382 189798 582326 190034
rect 582562 189798 582646 190034
rect 582882 189798 586302 190034
rect 586538 189798 586622 190034
rect 586858 189798 592650 190034
rect -8726 189766 592650 189798
rect -8726 185854 592650 185886
rect -8726 185618 -1974 185854
rect -1738 185618 -1654 185854
rect -1418 185618 5826 185854
rect 6062 185618 6146 185854
rect 6382 185618 185826 185854
rect 186062 185618 186146 185854
rect 186382 185618 221826 185854
rect 222062 185618 222146 185854
rect 222382 185618 257826 185854
rect 258062 185618 258146 185854
rect 258382 185618 293826 185854
rect 294062 185618 294146 185854
rect 294382 185618 329826 185854
rect 330062 185618 330146 185854
rect 330382 185618 365826 185854
rect 366062 185618 366146 185854
rect 366382 185618 401826 185854
rect 402062 185618 402146 185854
rect 402382 185618 570350 185854
rect 570586 185618 570670 185854
rect 570906 185618 585342 185854
rect 585578 185618 585662 185854
rect 585898 185618 592650 185854
rect -8726 185534 592650 185618
rect -8726 185298 -1974 185534
rect -1738 185298 -1654 185534
rect -1418 185298 5826 185534
rect 6062 185298 6146 185534
rect 6382 185298 185826 185534
rect 186062 185298 186146 185534
rect 186382 185298 221826 185534
rect 222062 185298 222146 185534
rect 222382 185298 257826 185534
rect 258062 185298 258146 185534
rect 258382 185298 293826 185534
rect 294062 185298 294146 185534
rect 294382 185298 329826 185534
rect 330062 185298 330146 185534
rect 330382 185298 365826 185534
rect 366062 185298 366146 185534
rect 366382 185298 401826 185534
rect 402062 185298 402146 185534
rect 402382 185298 570350 185534
rect 570586 185298 570670 185534
rect 570906 185298 585342 185534
rect 585578 185298 585662 185534
rect 585898 185298 592650 185534
rect -8726 185266 592650 185298
rect -8726 154354 592650 154386
rect -8726 154118 -2934 154354
rect -2698 154118 -2614 154354
rect -2378 154118 13198 154354
rect 13434 154118 13518 154354
rect 13754 154118 167826 154354
rect 168062 154118 168146 154354
rect 168382 154118 203826 154354
rect 204062 154118 204146 154354
rect 204382 154118 239826 154354
rect 240062 154118 240146 154354
rect 240382 154118 275826 154354
rect 276062 154118 276146 154354
rect 276382 154118 311826 154354
rect 312062 154118 312146 154354
rect 312382 154118 347826 154354
rect 348062 154118 348146 154354
rect 348382 154118 383826 154354
rect 384062 154118 384146 154354
rect 384382 154118 419826 154354
rect 420062 154118 420146 154354
rect 420382 154118 563826 154354
rect 564062 154118 564146 154354
rect 564382 154118 582326 154354
rect 582562 154118 582646 154354
rect 582882 154118 586302 154354
rect 586538 154118 586622 154354
rect 586858 154118 592650 154354
rect -8726 154034 592650 154118
rect -8726 153798 -2934 154034
rect -2698 153798 -2614 154034
rect -2378 153798 13198 154034
rect 13434 153798 13518 154034
rect 13754 153798 167826 154034
rect 168062 153798 168146 154034
rect 168382 153798 203826 154034
rect 204062 153798 204146 154034
rect 204382 153798 239826 154034
rect 240062 153798 240146 154034
rect 240382 153798 275826 154034
rect 276062 153798 276146 154034
rect 276382 153798 311826 154034
rect 312062 153798 312146 154034
rect 312382 153798 347826 154034
rect 348062 153798 348146 154034
rect 348382 153798 383826 154034
rect 384062 153798 384146 154034
rect 384382 153798 419826 154034
rect 420062 153798 420146 154034
rect 420382 153798 563826 154034
rect 564062 153798 564146 154034
rect 564382 153798 582326 154034
rect 582562 153798 582646 154034
rect 582882 153798 586302 154034
rect 586538 153798 586622 154034
rect 586858 153798 592650 154034
rect -8726 153766 592650 153798
rect -8726 149854 592650 149886
rect -8726 149618 -1974 149854
rect -1738 149618 -1654 149854
rect -1418 149618 5826 149854
rect 6062 149618 6146 149854
rect 6382 149618 185826 149854
rect 186062 149618 186146 149854
rect 186382 149618 221826 149854
rect 222062 149618 222146 149854
rect 222382 149618 257826 149854
rect 258062 149618 258146 149854
rect 258382 149618 293826 149854
rect 294062 149618 294146 149854
rect 294382 149618 329826 149854
rect 330062 149618 330146 149854
rect 330382 149618 365826 149854
rect 366062 149618 366146 149854
rect 366382 149618 401826 149854
rect 402062 149618 402146 149854
rect 402382 149618 570350 149854
rect 570586 149618 570670 149854
rect 570906 149618 585342 149854
rect 585578 149618 585662 149854
rect 585898 149618 592650 149854
rect -8726 149534 592650 149618
rect -8726 149298 -1974 149534
rect -1738 149298 -1654 149534
rect -1418 149298 5826 149534
rect 6062 149298 6146 149534
rect 6382 149298 185826 149534
rect 186062 149298 186146 149534
rect 186382 149298 221826 149534
rect 222062 149298 222146 149534
rect 222382 149298 257826 149534
rect 258062 149298 258146 149534
rect 258382 149298 293826 149534
rect 294062 149298 294146 149534
rect 294382 149298 329826 149534
rect 330062 149298 330146 149534
rect 330382 149298 365826 149534
rect 366062 149298 366146 149534
rect 366382 149298 401826 149534
rect 402062 149298 402146 149534
rect 402382 149298 570350 149534
rect 570586 149298 570670 149534
rect 570906 149298 585342 149534
rect 585578 149298 585662 149534
rect 585898 149298 592650 149534
rect -8726 149266 592650 149298
rect -8726 118354 592650 118386
rect -8726 118118 -2934 118354
rect -2698 118118 -2614 118354
rect -2378 118118 23826 118354
rect 24062 118118 24146 118354
rect 24382 118118 59826 118354
rect 60062 118118 60146 118354
rect 60382 118118 95826 118354
rect 96062 118118 96146 118354
rect 96382 118118 131826 118354
rect 132062 118118 132146 118354
rect 132382 118118 167826 118354
rect 168062 118118 168146 118354
rect 168382 118118 203826 118354
rect 204062 118118 204146 118354
rect 204382 118118 239826 118354
rect 240062 118118 240146 118354
rect 240382 118118 275826 118354
rect 276062 118118 276146 118354
rect 276382 118118 311826 118354
rect 312062 118118 312146 118354
rect 312382 118118 347826 118354
rect 348062 118118 348146 118354
rect 348382 118118 383826 118354
rect 384062 118118 384146 118354
rect 384382 118118 419826 118354
rect 420062 118118 420146 118354
rect 420382 118118 455826 118354
rect 456062 118118 456146 118354
rect 456382 118118 491826 118354
rect 492062 118118 492146 118354
rect 492382 118118 527826 118354
rect 528062 118118 528146 118354
rect 528382 118118 563826 118354
rect 564062 118118 564146 118354
rect 564382 118118 582326 118354
rect 582562 118118 582646 118354
rect 582882 118118 586302 118354
rect 586538 118118 586622 118354
rect 586858 118118 592650 118354
rect -8726 118034 592650 118118
rect -8726 117798 -2934 118034
rect -2698 117798 -2614 118034
rect -2378 117798 23826 118034
rect 24062 117798 24146 118034
rect 24382 117798 59826 118034
rect 60062 117798 60146 118034
rect 60382 117798 95826 118034
rect 96062 117798 96146 118034
rect 96382 117798 131826 118034
rect 132062 117798 132146 118034
rect 132382 117798 167826 118034
rect 168062 117798 168146 118034
rect 168382 117798 203826 118034
rect 204062 117798 204146 118034
rect 204382 117798 239826 118034
rect 240062 117798 240146 118034
rect 240382 117798 275826 118034
rect 276062 117798 276146 118034
rect 276382 117798 311826 118034
rect 312062 117798 312146 118034
rect 312382 117798 347826 118034
rect 348062 117798 348146 118034
rect 348382 117798 383826 118034
rect 384062 117798 384146 118034
rect 384382 117798 419826 118034
rect 420062 117798 420146 118034
rect 420382 117798 455826 118034
rect 456062 117798 456146 118034
rect 456382 117798 491826 118034
rect 492062 117798 492146 118034
rect 492382 117798 527826 118034
rect 528062 117798 528146 118034
rect 528382 117798 563826 118034
rect 564062 117798 564146 118034
rect 564382 117798 582326 118034
rect 582562 117798 582646 118034
rect 582882 117798 586302 118034
rect 586538 117798 586622 118034
rect 586858 117798 592650 118034
rect -8726 117766 592650 117798
rect -8726 113854 592650 113886
rect -8726 113618 -1974 113854
rect -1738 113618 -1654 113854
rect -1418 113618 5826 113854
rect 6062 113618 6146 113854
rect 6382 113715 293826 113854
rect 6382 113618 41826 113715
rect -8726 113534 41826 113618
rect -8726 113298 -1974 113534
rect -1738 113298 -1654 113534
rect -1418 113298 5826 113534
rect 6062 113298 6146 113534
rect 6382 113479 41826 113534
rect 42062 113479 42146 113715
rect 42382 113479 77826 113715
rect 78062 113479 78146 113715
rect 78382 113479 113826 113715
rect 114062 113479 114146 113715
rect 114382 113479 149826 113715
rect 150062 113479 150146 113715
rect 150382 113618 293826 113715
rect 294062 113618 294146 113854
rect 294382 113618 401826 113854
rect 402062 113618 402146 113854
rect 402382 113715 585342 113854
rect 402382 113618 437826 113715
rect 150382 113534 437826 113618
rect 150382 113479 293826 113534
rect 6382 113298 293826 113479
rect 294062 113298 294146 113534
rect 294382 113298 401826 113534
rect 402062 113298 402146 113534
rect 402382 113479 437826 113534
rect 438062 113479 438146 113715
rect 438382 113479 473826 113715
rect 474062 113479 474146 113715
rect 474382 113479 509826 113715
rect 510062 113479 510146 113715
rect 510382 113479 545826 113715
rect 546062 113479 546146 113715
rect 546382 113618 585342 113715
rect 585578 113618 585662 113854
rect 585898 113618 592650 113854
rect 546382 113534 592650 113618
rect 546382 113479 585342 113534
rect 402382 113298 585342 113479
rect 585578 113298 585662 113534
rect 585898 113298 592650 113534
rect -8726 113266 592650 113298
rect -8726 82354 592650 82386
rect -8726 82118 -2934 82354
rect -2698 82118 -2614 82354
rect -2378 82118 13198 82354
rect 13434 82118 13518 82354
rect 13754 82118 167826 82354
rect 168062 82118 168146 82354
rect 168382 82118 291590 82354
rect 291826 82118 291910 82354
rect 292146 82118 419826 82354
rect 420062 82118 420146 82354
rect 420382 82118 563826 82354
rect 564062 82118 564146 82354
rect 564382 82118 582326 82354
rect 582562 82118 582646 82354
rect 582882 82118 586302 82354
rect 586538 82118 586622 82354
rect 586858 82118 592650 82354
rect -8726 82034 592650 82118
rect -8726 81798 -2934 82034
rect -2698 81798 -2614 82034
rect -2378 81798 13198 82034
rect 13434 81798 13518 82034
rect 13754 81798 167826 82034
rect 168062 81798 168146 82034
rect 168382 81798 291590 82034
rect 291826 81798 291910 82034
rect 292146 81798 419826 82034
rect 420062 81798 420146 82034
rect 420382 81798 563826 82034
rect 564062 81798 564146 82034
rect 564382 81798 582326 82034
rect 582562 81798 582646 82034
rect 582882 81798 586302 82034
rect 586538 81798 586622 82034
rect 586858 81798 592650 82034
rect -8726 81766 592650 81798
rect -8726 77854 592650 77886
rect -8726 77618 -1974 77854
rect -1738 77618 -1654 77854
rect -1418 77618 5826 77854
rect 6062 77618 6146 77854
rect 6382 77618 173094 77854
rect 173330 77618 173414 77854
rect 173650 77618 293826 77854
rect 294062 77618 294146 77854
rect 294382 77618 401826 77854
rect 402062 77618 402146 77854
rect 402382 77618 570350 77854
rect 570586 77618 570670 77854
rect 570906 77618 585342 77854
rect 585578 77618 585662 77854
rect 585898 77618 592650 77854
rect -8726 77534 592650 77618
rect -8726 77298 -1974 77534
rect -1738 77298 -1654 77534
rect -1418 77298 5826 77534
rect 6062 77298 6146 77534
rect 6382 77298 173094 77534
rect 173330 77298 173414 77534
rect 173650 77298 293826 77534
rect 294062 77298 294146 77534
rect 294382 77298 401826 77534
rect 402062 77298 402146 77534
rect 402382 77298 570350 77534
rect 570586 77298 570670 77534
rect 570906 77298 585342 77534
rect 585578 77298 585662 77534
rect 585898 77298 592650 77534
rect -8726 77266 592650 77298
rect -8726 46354 592650 46386
rect -8726 46118 -2934 46354
rect -2698 46118 -2614 46354
rect -2378 46118 13198 46354
rect 13434 46118 13518 46354
rect 13754 46118 167826 46354
rect 168062 46118 168146 46354
rect 168382 46118 291590 46354
rect 291826 46118 291910 46354
rect 292146 46118 419826 46354
rect 420062 46118 420146 46354
rect 420382 46118 563826 46354
rect 564062 46118 564146 46354
rect 564382 46118 582326 46354
rect 582562 46118 582646 46354
rect 582882 46118 586302 46354
rect 586538 46118 586622 46354
rect 586858 46118 592650 46354
rect -8726 46034 592650 46118
rect -8726 45798 -2934 46034
rect -2698 45798 -2614 46034
rect -2378 45798 13198 46034
rect 13434 45798 13518 46034
rect 13754 45798 167826 46034
rect 168062 45798 168146 46034
rect 168382 45798 291590 46034
rect 291826 45798 291910 46034
rect 292146 45798 419826 46034
rect 420062 45798 420146 46034
rect 420382 45798 563826 46034
rect 564062 45798 564146 46034
rect 564382 45798 582326 46034
rect 582562 45798 582646 46034
rect 582882 45798 586302 46034
rect 586538 45798 586622 46034
rect 586858 45798 592650 46034
rect -8726 45766 592650 45798
rect -8726 41854 592650 41886
rect -8726 41618 -1974 41854
rect -1738 41618 -1654 41854
rect -1418 41618 5826 41854
rect 6062 41618 6146 41854
rect 6382 41618 173094 41854
rect 173330 41618 173414 41854
rect 173650 41618 293826 41854
rect 294062 41618 294146 41854
rect 294382 41618 401826 41854
rect 402062 41618 402146 41854
rect 402382 41618 570350 41854
rect 570586 41618 570670 41854
rect 570906 41618 585342 41854
rect 585578 41618 585662 41854
rect 585898 41618 592650 41854
rect -8726 41534 592650 41618
rect -8726 41298 -1974 41534
rect -1738 41298 -1654 41534
rect -1418 41298 5826 41534
rect 6062 41298 6146 41534
rect 6382 41298 173094 41534
rect 173330 41298 173414 41534
rect 173650 41298 293826 41534
rect 294062 41298 294146 41534
rect 294382 41298 401826 41534
rect 402062 41298 402146 41534
rect 402382 41298 570350 41534
rect 570586 41298 570670 41534
rect 570906 41298 585342 41534
rect 585578 41298 585662 41534
rect 585898 41298 592650 41534
rect -8726 41266 592650 41298
rect -8726 10354 592650 10386
rect -8726 10118 -2934 10354
rect -2698 10118 -2614 10354
rect -2378 10118 23826 10354
rect 24062 10118 24146 10354
rect 24382 10118 59826 10354
rect 60062 10118 60146 10354
rect 60382 10118 95826 10354
rect 96062 10118 96146 10354
rect 96382 10118 131826 10354
rect 132062 10118 132146 10354
rect 132382 10118 167826 10354
rect 168062 10118 168146 10354
rect 168382 10118 203826 10354
rect 204062 10118 204146 10354
rect 204382 10118 239826 10354
rect 240062 10118 240146 10354
rect 240382 10118 275826 10354
rect 276062 10118 276146 10354
rect 276382 10118 311826 10354
rect 312062 10118 312146 10354
rect 312382 10118 347826 10354
rect 348062 10118 348146 10354
rect 348382 10118 383826 10354
rect 384062 10118 384146 10354
rect 384382 10118 419826 10354
rect 420062 10118 420146 10354
rect 420382 10118 455826 10354
rect 456062 10118 456146 10354
rect 456382 10118 491826 10354
rect 492062 10118 492146 10354
rect 492382 10118 527826 10354
rect 528062 10118 528146 10354
rect 528382 10118 563826 10354
rect 564062 10118 564146 10354
rect 564382 10118 582326 10354
rect 582562 10118 582646 10354
rect 582882 10118 586302 10354
rect 586538 10118 586622 10354
rect 586858 10118 592650 10354
rect -8726 10034 592650 10118
rect -8726 9798 -2934 10034
rect -2698 9798 -2614 10034
rect -2378 9798 23826 10034
rect 24062 9798 24146 10034
rect 24382 9798 59826 10034
rect 60062 9798 60146 10034
rect 60382 9798 95826 10034
rect 96062 9798 96146 10034
rect 96382 9798 131826 10034
rect 132062 9798 132146 10034
rect 132382 9798 167826 10034
rect 168062 9798 168146 10034
rect 168382 9798 203826 10034
rect 204062 9798 204146 10034
rect 204382 9798 239826 10034
rect 240062 9798 240146 10034
rect 240382 9798 275826 10034
rect 276062 9798 276146 10034
rect 276382 9798 311826 10034
rect 312062 9798 312146 10034
rect 312382 9798 347826 10034
rect 348062 9798 348146 10034
rect 348382 9798 383826 10034
rect 384062 9798 384146 10034
rect 384382 9798 419826 10034
rect 420062 9798 420146 10034
rect 420382 9798 455826 10034
rect 456062 9798 456146 10034
rect 456382 9798 491826 10034
rect 492062 9798 492146 10034
rect 492382 9798 527826 10034
rect 528062 9798 528146 10034
rect 528382 9798 563826 10034
rect 564062 9798 564146 10034
rect 564382 9798 582326 10034
rect 582562 9798 582646 10034
rect 582882 9798 586302 10034
rect 586538 9798 586622 10034
rect 586858 9798 592650 10034
rect -8726 9766 592650 9798
rect -8726 5854 592650 5886
rect -8726 5618 -1974 5854
rect -1738 5618 -1654 5854
rect -1418 5618 585342 5854
rect 585578 5618 585662 5854
rect 585898 5618 592650 5854
rect -8726 5534 592650 5618
rect -8726 5298 -1974 5534
rect -1738 5298 -1654 5534
rect -1418 5298 585342 5534
rect 585578 5298 585662 5534
rect 585898 5298 592650 5534
rect -8726 5266 592650 5298
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 582326 -1306
rect 582562 -1542 582646 -1306
rect 582882 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 582326 -1626
rect 582562 -1862 582646 -1626
rect 582882 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use Marmot  Marmot
timestamp 0
transform 1 0 4000 0 1 4000
box -960 -960 576960 696960
<< labels >>
flabel metal3 s 583520 285276 584960 285516 0 FreeSans 960 0 0 0 analog_io[0]
port 0 nsew signal bidirectional
flabel metal2 s 446098 703520 446210 704960 0 FreeSans 448 90 0 0 analog_io[10]
port 1 nsew signal bidirectional
flabel metal2 s 381146 703520 381258 704960 0 FreeSans 448 90 0 0 analog_io[11]
port 2 nsew signal bidirectional
flabel metal2 s 316286 703520 316398 704960 0 FreeSans 448 90 0 0 analog_io[12]
port 3 nsew signal bidirectional
flabel metal2 s 251426 703520 251538 704960 0 FreeSans 448 90 0 0 analog_io[13]
port 4 nsew signal bidirectional
flabel metal2 s 186474 703520 186586 704960 0 FreeSans 448 90 0 0 analog_io[14]
port 5 nsew signal bidirectional
flabel metal2 s 121614 703520 121726 704960 0 FreeSans 448 90 0 0 analog_io[15]
port 6 nsew signal bidirectional
flabel metal2 s 56754 703520 56866 704960 0 FreeSans 448 90 0 0 analog_io[16]
port 7 nsew signal bidirectional
flabel metal3 s -960 697220 480 697460 0 FreeSans 960 0 0 0 analog_io[17]
port 8 nsew signal bidirectional
flabel metal3 s -960 644996 480 645236 0 FreeSans 960 0 0 0 analog_io[18]
port 9 nsew signal bidirectional
flabel metal3 s -960 592908 480 593148 0 FreeSans 960 0 0 0 analog_io[19]
port 10 nsew signal bidirectional
flabel metal3 s 583520 338452 584960 338692 0 FreeSans 960 0 0 0 analog_io[1]
port 11 nsew signal bidirectional
flabel metal3 s -960 540684 480 540924 0 FreeSans 960 0 0 0 analog_io[20]
port 12 nsew signal bidirectional
flabel metal3 s -960 488596 480 488836 0 FreeSans 960 0 0 0 analog_io[21]
port 13 nsew signal bidirectional
flabel metal3 s -960 436508 480 436748 0 FreeSans 960 0 0 0 analog_io[22]
port 14 nsew signal bidirectional
flabel metal3 s -960 384284 480 384524 0 FreeSans 960 0 0 0 analog_io[23]
port 15 nsew signal bidirectional
flabel metal3 s -960 332196 480 332436 0 FreeSans 960 0 0 0 analog_io[24]
port 16 nsew signal bidirectional
flabel metal3 s -960 279972 480 280212 0 FreeSans 960 0 0 0 analog_io[25]
port 17 nsew signal bidirectional
flabel metal3 s -960 227884 480 228124 0 FreeSans 960 0 0 0 analog_io[26]
port 18 nsew signal bidirectional
flabel metal3 s -960 175796 480 176036 0 FreeSans 960 0 0 0 analog_io[27]
port 19 nsew signal bidirectional
flabel metal3 s -960 123572 480 123812 0 FreeSans 960 0 0 0 analog_io[28]
port 20 nsew signal bidirectional
flabel metal3 s 583520 391628 584960 391868 0 FreeSans 960 0 0 0 analog_io[2]
port 21 nsew signal bidirectional
flabel metal3 s 583520 444668 584960 444908 0 FreeSans 960 0 0 0 analog_io[3]
port 22 nsew signal bidirectional
flabel metal3 s 583520 497844 584960 498084 0 FreeSans 960 0 0 0 analog_io[4]
port 23 nsew signal bidirectional
flabel metal3 s 583520 551020 584960 551260 0 FreeSans 960 0 0 0 analog_io[5]
port 24 nsew signal bidirectional
flabel metal3 s 583520 604060 584960 604300 0 FreeSans 960 0 0 0 analog_io[6]
port 25 nsew signal bidirectional
flabel metal3 s 583520 657236 584960 657476 0 FreeSans 960 0 0 0 analog_io[7]
port 26 nsew signal bidirectional
flabel metal2 s 575818 703520 575930 704960 0 FreeSans 448 90 0 0 analog_io[8]
port 27 nsew signal bidirectional
flabel metal2 s 510958 703520 511070 704960 0 FreeSans 448 90 0 0 analog_io[9]
port 28 nsew signal bidirectional
flabel metal3 s 583520 6476 584960 6716 0 FreeSans 960 0 0 0 io_in[0]
port 29 nsew signal input
flabel metal3 s 583520 457996 584960 458236 0 FreeSans 960 0 0 0 io_in[10]
port 30 nsew signal input
flabel metal3 s 583520 511172 584960 511412 0 FreeSans 960 0 0 0 io_in[11]
port 31 nsew signal input
flabel metal3 s 583520 564212 584960 564452 0 FreeSans 960 0 0 0 io_in[12]
port 32 nsew signal input
flabel metal3 s 583520 617388 584960 617628 0 FreeSans 960 0 0 0 io_in[13]
port 33 nsew signal input
flabel metal3 s 583520 670564 584960 670804 0 FreeSans 960 0 0 0 io_in[14]
port 34 nsew signal input
flabel metal2 s 559626 703520 559738 704960 0 FreeSans 448 90 0 0 io_in[15]
port 35 nsew signal input
flabel metal2 s 494766 703520 494878 704960 0 FreeSans 448 90 0 0 io_in[16]
port 36 nsew signal input
flabel metal2 s 429814 703520 429926 704960 0 FreeSans 448 90 0 0 io_in[17]
port 37 nsew signal input
flabel metal2 s 364954 703520 365066 704960 0 FreeSans 448 90 0 0 io_in[18]
port 38 nsew signal input
flabel metal2 s 300094 703520 300206 704960 0 FreeSans 448 90 0 0 io_in[19]
port 39 nsew signal input
flabel metal3 s 583520 46188 584960 46428 0 FreeSans 960 0 0 0 io_in[1]
port 40 nsew signal input
flabel metal2 s 235142 703520 235254 704960 0 FreeSans 448 90 0 0 io_in[20]
port 41 nsew signal input
flabel metal2 s 170282 703520 170394 704960 0 FreeSans 448 90 0 0 io_in[21]
port 42 nsew signal input
flabel metal2 s 105422 703520 105534 704960 0 FreeSans 448 90 0 0 io_in[22]
port 43 nsew signal input
flabel metal2 s 40470 703520 40582 704960 0 FreeSans 448 90 0 0 io_in[23]
port 44 nsew signal input
flabel metal3 s -960 684164 480 684404 0 FreeSans 960 0 0 0 io_in[24]
port 45 nsew signal input
flabel metal3 s -960 631940 480 632180 0 FreeSans 960 0 0 0 io_in[25]
port 46 nsew signal input
flabel metal3 s -960 579852 480 580092 0 FreeSans 960 0 0 0 io_in[26]
port 47 nsew signal input
flabel metal3 s -960 527764 480 528004 0 FreeSans 960 0 0 0 io_in[27]
port 48 nsew signal input
flabel metal3 s -960 475540 480 475780 0 FreeSans 960 0 0 0 io_in[28]
port 49 nsew signal input
flabel metal3 s -960 423452 480 423692 0 FreeSans 960 0 0 0 io_in[29]
port 50 nsew signal input
flabel metal3 s 583520 86036 584960 86276 0 FreeSans 960 0 0 0 io_in[2]
port 51 nsew signal input
flabel metal3 s -960 371228 480 371468 0 FreeSans 960 0 0 0 io_in[30]
port 52 nsew signal input
flabel metal3 s -960 319140 480 319380 0 FreeSans 960 0 0 0 io_in[31]
port 53 nsew signal input
flabel metal3 s -960 267052 480 267292 0 FreeSans 960 0 0 0 io_in[32]
port 54 nsew signal input
flabel metal3 s -960 214828 480 215068 0 FreeSans 960 0 0 0 io_in[33]
port 55 nsew signal input
flabel metal3 s -960 162740 480 162980 0 FreeSans 960 0 0 0 io_in[34]
port 56 nsew signal input
flabel metal3 s -960 110516 480 110756 0 FreeSans 960 0 0 0 io_in[35]
port 57 nsew signal input
flabel metal3 s -960 71484 480 71724 0 FreeSans 960 0 0 0 io_in[36]
port 58 nsew signal input
flabel metal3 s -960 32316 480 32556 0 FreeSans 960 0 0 0 io_in[37]
port 59 nsew signal input
flabel metal3 s 583520 125884 584960 126124 0 FreeSans 960 0 0 0 io_in[3]
port 60 nsew signal input
flabel metal3 s 583520 165732 584960 165972 0 FreeSans 960 0 0 0 io_in[4]
port 61 nsew signal input
flabel metal3 s 583520 205580 584960 205820 0 FreeSans 960 0 0 0 io_in[5]
port 62 nsew signal input
flabel metal3 s 583520 245428 584960 245668 0 FreeSans 960 0 0 0 io_in[6]
port 63 nsew signal input
flabel metal3 s 583520 298604 584960 298844 0 FreeSans 960 0 0 0 io_in[7]
port 64 nsew signal input
flabel metal3 s 583520 351780 584960 352020 0 FreeSans 960 0 0 0 io_in[8]
port 65 nsew signal input
flabel metal3 s 583520 404820 584960 405060 0 FreeSans 960 0 0 0 io_in[9]
port 66 nsew signal input
flabel metal3 s 583520 32996 584960 33236 0 FreeSans 960 0 0 0 io_oeb[0]
port 67 nsew signal tristate
flabel metal3 s 583520 484516 584960 484756 0 FreeSans 960 0 0 0 io_oeb[10]
port 68 nsew signal tristate
flabel metal3 s 583520 537692 584960 537932 0 FreeSans 960 0 0 0 io_oeb[11]
port 69 nsew signal tristate
flabel metal3 s 583520 590868 584960 591108 0 FreeSans 960 0 0 0 io_oeb[12]
port 70 nsew signal tristate
flabel metal3 s 583520 643908 584960 644148 0 FreeSans 960 0 0 0 io_oeb[13]
port 71 nsew signal tristate
flabel metal3 s 583520 697084 584960 697324 0 FreeSans 960 0 0 0 io_oeb[14]
port 72 nsew signal tristate
flabel metal2 s 527150 703520 527262 704960 0 FreeSans 448 90 0 0 io_oeb[15]
port 73 nsew signal tristate
flabel metal2 s 462290 703520 462402 704960 0 FreeSans 448 90 0 0 io_oeb[16]
port 74 nsew signal tristate
flabel metal2 s 397430 703520 397542 704960 0 FreeSans 448 90 0 0 io_oeb[17]
port 75 nsew signal tristate
flabel metal2 s 332478 703520 332590 704960 0 FreeSans 448 90 0 0 io_oeb[18]
port 76 nsew signal tristate
flabel metal2 s 267618 703520 267730 704960 0 FreeSans 448 90 0 0 io_oeb[19]
port 77 nsew signal tristate
flabel metal3 s 583520 72844 584960 73084 0 FreeSans 960 0 0 0 io_oeb[1]
port 78 nsew signal tristate
flabel metal2 s 202758 703520 202870 704960 0 FreeSans 448 90 0 0 io_oeb[20]
port 79 nsew signal tristate
flabel metal2 s 137806 703520 137918 704960 0 FreeSans 448 90 0 0 io_oeb[21]
port 80 nsew signal tristate
flabel metal2 s 72946 703520 73058 704960 0 FreeSans 448 90 0 0 io_oeb[22]
port 81 nsew signal tristate
flabel metal2 s 8086 703520 8198 704960 0 FreeSans 448 90 0 0 io_oeb[23]
port 82 nsew signal tristate
flabel metal3 s -960 658052 480 658292 0 FreeSans 960 0 0 0 io_oeb[24]
port 83 nsew signal tristate
flabel metal3 s -960 605964 480 606204 0 FreeSans 960 0 0 0 io_oeb[25]
port 84 nsew signal tristate
flabel metal3 s -960 553740 480 553980 0 FreeSans 960 0 0 0 io_oeb[26]
port 85 nsew signal tristate
flabel metal3 s -960 501652 480 501892 0 FreeSans 960 0 0 0 io_oeb[27]
port 86 nsew signal tristate
flabel metal3 s -960 449428 480 449668 0 FreeSans 960 0 0 0 io_oeb[28]
port 87 nsew signal tristate
flabel metal3 s -960 397340 480 397580 0 FreeSans 960 0 0 0 io_oeb[29]
port 88 nsew signal tristate
flabel metal3 s 583520 112692 584960 112932 0 FreeSans 960 0 0 0 io_oeb[2]
port 89 nsew signal tristate
flabel metal3 s -960 345252 480 345492 0 FreeSans 960 0 0 0 io_oeb[30]
port 90 nsew signal tristate
flabel metal3 s -960 293028 480 293268 0 FreeSans 960 0 0 0 io_oeb[31]
port 91 nsew signal tristate
flabel metal3 s -960 240940 480 241180 0 FreeSans 960 0 0 0 io_oeb[32]
port 92 nsew signal tristate
flabel metal3 s -960 188716 480 188956 0 FreeSans 960 0 0 0 io_oeb[33]
port 93 nsew signal tristate
flabel metal3 s -960 136628 480 136868 0 FreeSans 960 0 0 0 io_oeb[34]
port 94 nsew signal tristate
flabel metal3 s -960 84540 480 84780 0 FreeSans 960 0 0 0 io_oeb[35]
port 95 nsew signal tristate
flabel metal3 s -960 45372 480 45612 0 FreeSans 960 0 0 0 io_oeb[36]
port 96 nsew signal tristate
flabel metal3 s -960 6340 480 6580 0 FreeSans 960 0 0 0 io_oeb[37]
port 97 nsew signal tristate
flabel metal3 s 583520 152540 584960 152780 0 FreeSans 960 0 0 0 io_oeb[3]
port 98 nsew signal tristate
flabel metal3 s 583520 192388 584960 192628 0 FreeSans 960 0 0 0 io_oeb[4]
port 99 nsew signal tristate
flabel metal3 s 583520 232236 584960 232476 0 FreeSans 960 0 0 0 io_oeb[5]
port 100 nsew signal tristate
flabel metal3 s 583520 272084 584960 272324 0 FreeSans 960 0 0 0 io_oeb[6]
port 101 nsew signal tristate
flabel metal3 s 583520 325124 584960 325364 0 FreeSans 960 0 0 0 io_oeb[7]
port 102 nsew signal tristate
flabel metal3 s 583520 378300 584960 378540 0 FreeSans 960 0 0 0 io_oeb[8]
port 103 nsew signal tristate
flabel metal3 s 583520 431476 584960 431716 0 FreeSans 960 0 0 0 io_oeb[9]
port 104 nsew signal tristate
flabel metal3 s 583520 19668 584960 19908 0 FreeSans 960 0 0 0 io_out[0]
port 105 nsew signal tristate
flabel metal3 s 583520 471324 584960 471564 0 FreeSans 960 0 0 0 io_out[10]
port 106 nsew signal tristate
flabel metal3 s 583520 524364 584960 524604 0 FreeSans 960 0 0 0 io_out[11]
port 107 nsew signal tristate
flabel metal3 s 583520 577540 584960 577780 0 FreeSans 960 0 0 0 io_out[12]
port 108 nsew signal tristate
flabel metal3 s 583520 630716 584960 630956 0 FreeSans 960 0 0 0 io_out[13]
port 109 nsew signal tristate
flabel metal3 s 583520 683756 584960 683996 0 FreeSans 960 0 0 0 io_out[14]
port 110 nsew signal tristate
flabel metal2 s 543434 703520 543546 704960 0 FreeSans 448 90 0 0 io_out[15]
port 111 nsew signal tristate
flabel metal2 s 478482 703520 478594 704960 0 FreeSans 448 90 0 0 io_out[16]
port 112 nsew signal tristate
flabel metal2 s 413622 703520 413734 704960 0 FreeSans 448 90 0 0 io_out[17]
port 113 nsew signal tristate
flabel metal2 s 348762 703520 348874 704960 0 FreeSans 448 90 0 0 io_out[18]
port 114 nsew signal tristate
flabel metal2 s 283810 703520 283922 704960 0 FreeSans 448 90 0 0 io_out[19]
port 115 nsew signal tristate
flabel metal3 s 583520 59516 584960 59756 0 FreeSans 960 0 0 0 io_out[1]
port 116 nsew signal tristate
flabel metal2 s 218950 703520 219062 704960 0 FreeSans 448 90 0 0 io_out[20]
port 117 nsew signal tristate
flabel metal2 s 154090 703520 154202 704960 0 FreeSans 448 90 0 0 io_out[21]
port 118 nsew signal tristate
flabel metal2 s 89138 703520 89250 704960 0 FreeSans 448 90 0 0 io_out[22]
port 119 nsew signal tristate
flabel metal2 s 24278 703520 24390 704960 0 FreeSans 448 90 0 0 io_out[23]
port 120 nsew signal tristate
flabel metal3 s -960 671108 480 671348 0 FreeSans 960 0 0 0 io_out[24]
port 121 nsew signal tristate
flabel metal3 s -960 619020 480 619260 0 FreeSans 960 0 0 0 io_out[25]
port 122 nsew signal tristate
flabel metal3 s -960 566796 480 567036 0 FreeSans 960 0 0 0 io_out[26]
port 123 nsew signal tristate
flabel metal3 s -960 514708 480 514948 0 FreeSans 960 0 0 0 io_out[27]
port 124 nsew signal tristate
flabel metal3 s -960 462484 480 462724 0 FreeSans 960 0 0 0 io_out[28]
port 125 nsew signal tristate
flabel metal3 s -960 410396 480 410636 0 FreeSans 960 0 0 0 io_out[29]
port 126 nsew signal tristate
flabel metal3 s 583520 99364 584960 99604 0 FreeSans 960 0 0 0 io_out[2]
port 127 nsew signal tristate
flabel metal3 s -960 358308 480 358548 0 FreeSans 960 0 0 0 io_out[30]
port 128 nsew signal tristate
flabel metal3 s -960 306084 480 306324 0 FreeSans 960 0 0 0 io_out[31]
port 129 nsew signal tristate
flabel metal3 s -960 253996 480 254236 0 FreeSans 960 0 0 0 io_out[32]
port 130 nsew signal tristate
flabel metal3 s -960 201772 480 202012 0 FreeSans 960 0 0 0 io_out[33]
port 131 nsew signal tristate
flabel metal3 s -960 149684 480 149924 0 FreeSans 960 0 0 0 io_out[34]
port 132 nsew signal tristate
flabel metal3 s -960 97460 480 97700 0 FreeSans 960 0 0 0 io_out[35]
port 133 nsew signal tristate
flabel metal3 s -960 58428 480 58668 0 FreeSans 960 0 0 0 io_out[36]
port 134 nsew signal tristate
flabel metal3 s -960 19260 480 19500 0 FreeSans 960 0 0 0 io_out[37]
port 135 nsew signal tristate
flabel metal3 s 583520 139212 584960 139452 0 FreeSans 960 0 0 0 io_out[3]
port 136 nsew signal tristate
flabel metal3 s 583520 179060 584960 179300 0 FreeSans 960 0 0 0 io_out[4]
port 137 nsew signal tristate
flabel metal3 s 583520 218908 584960 219148 0 FreeSans 960 0 0 0 io_out[5]
port 138 nsew signal tristate
flabel metal3 s 583520 258756 584960 258996 0 FreeSans 960 0 0 0 io_out[6]
port 139 nsew signal tristate
flabel metal3 s 583520 311932 584960 312172 0 FreeSans 960 0 0 0 io_out[7]
port 140 nsew signal tristate
flabel metal3 s 583520 364972 584960 365212 0 FreeSans 960 0 0 0 io_out[8]
port 141 nsew signal tristate
flabel metal3 s 583520 418148 584960 418388 0 FreeSans 960 0 0 0 io_out[9]
port 142 nsew signal tristate
flabel metal2 s 125846 -960 125958 480 0 FreeSans 448 90 0 0 la_data_in[0]
port 143 nsew signal input
flabel metal2 s 480506 -960 480618 480 0 FreeSans 448 90 0 0 la_data_in[100]
port 144 nsew signal input
flabel metal2 s 484002 -960 484114 480 0 FreeSans 448 90 0 0 la_data_in[101]
port 145 nsew signal input
flabel metal2 s 487590 -960 487702 480 0 FreeSans 448 90 0 0 la_data_in[102]
port 146 nsew signal input
flabel metal2 s 491086 -960 491198 480 0 FreeSans 448 90 0 0 la_data_in[103]
port 147 nsew signal input
flabel metal2 s 494674 -960 494786 480 0 FreeSans 448 90 0 0 la_data_in[104]
port 148 nsew signal input
flabel metal2 s 498170 -960 498282 480 0 FreeSans 448 90 0 0 la_data_in[105]
port 149 nsew signal input
flabel metal2 s 501758 -960 501870 480 0 FreeSans 448 90 0 0 la_data_in[106]
port 150 nsew signal input
flabel metal2 s 505346 -960 505458 480 0 FreeSans 448 90 0 0 la_data_in[107]
port 151 nsew signal input
flabel metal2 s 508842 -960 508954 480 0 FreeSans 448 90 0 0 la_data_in[108]
port 152 nsew signal input
flabel metal2 s 512430 -960 512542 480 0 FreeSans 448 90 0 0 la_data_in[109]
port 153 nsew signal input
flabel metal2 s 161266 -960 161378 480 0 FreeSans 448 90 0 0 la_data_in[10]
port 154 nsew signal input
flabel metal2 s 515926 -960 516038 480 0 FreeSans 448 90 0 0 la_data_in[110]
port 155 nsew signal input
flabel metal2 s 519514 -960 519626 480 0 FreeSans 448 90 0 0 la_data_in[111]
port 156 nsew signal input
flabel metal2 s 523010 -960 523122 480 0 FreeSans 448 90 0 0 la_data_in[112]
port 157 nsew signal input
flabel metal2 s 526598 -960 526710 480 0 FreeSans 448 90 0 0 la_data_in[113]
port 158 nsew signal input
flabel metal2 s 530094 -960 530206 480 0 FreeSans 448 90 0 0 la_data_in[114]
port 159 nsew signal input
flabel metal2 s 533682 -960 533794 480 0 FreeSans 448 90 0 0 la_data_in[115]
port 160 nsew signal input
flabel metal2 s 537178 -960 537290 480 0 FreeSans 448 90 0 0 la_data_in[116]
port 161 nsew signal input
flabel metal2 s 540766 -960 540878 480 0 FreeSans 448 90 0 0 la_data_in[117]
port 162 nsew signal input
flabel metal2 s 544354 -960 544466 480 0 FreeSans 448 90 0 0 la_data_in[118]
port 163 nsew signal input
flabel metal2 s 547850 -960 547962 480 0 FreeSans 448 90 0 0 la_data_in[119]
port 164 nsew signal input
flabel metal2 s 164854 -960 164966 480 0 FreeSans 448 90 0 0 la_data_in[11]
port 165 nsew signal input
flabel metal2 s 551438 -960 551550 480 0 FreeSans 448 90 0 0 la_data_in[120]
port 166 nsew signal input
flabel metal2 s 554934 -960 555046 480 0 FreeSans 448 90 0 0 la_data_in[121]
port 167 nsew signal input
flabel metal2 s 558522 -960 558634 480 0 FreeSans 448 90 0 0 la_data_in[122]
port 168 nsew signal input
flabel metal2 s 562018 -960 562130 480 0 FreeSans 448 90 0 0 la_data_in[123]
port 169 nsew signal input
flabel metal2 s 565606 -960 565718 480 0 FreeSans 448 90 0 0 la_data_in[124]
port 170 nsew signal input
flabel metal2 s 569102 -960 569214 480 0 FreeSans 448 90 0 0 la_data_in[125]
port 171 nsew signal input
flabel metal2 s 572690 -960 572802 480 0 FreeSans 448 90 0 0 la_data_in[126]
port 172 nsew signal input
flabel metal2 s 576278 -960 576390 480 0 FreeSans 448 90 0 0 la_data_in[127]
port 173 nsew signal input
flabel metal2 s 168350 -960 168462 480 0 FreeSans 448 90 0 0 la_data_in[12]
port 174 nsew signal input
flabel metal2 s 171938 -960 172050 480 0 FreeSans 448 90 0 0 la_data_in[13]
port 175 nsew signal input
flabel metal2 s 175434 -960 175546 480 0 FreeSans 448 90 0 0 la_data_in[14]
port 176 nsew signal input
flabel metal2 s 179022 -960 179134 480 0 FreeSans 448 90 0 0 la_data_in[15]
port 177 nsew signal input
flabel metal2 s 182518 -960 182630 480 0 FreeSans 448 90 0 0 la_data_in[16]
port 178 nsew signal input
flabel metal2 s 186106 -960 186218 480 0 FreeSans 448 90 0 0 la_data_in[17]
port 179 nsew signal input
flabel metal2 s 189694 -960 189806 480 0 FreeSans 448 90 0 0 la_data_in[18]
port 180 nsew signal input
flabel metal2 s 193190 -960 193302 480 0 FreeSans 448 90 0 0 la_data_in[19]
port 181 nsew signal input
flabel metal2 s 129342 -960 129454 480 0 FreeSans 448 90 0 0 la_data_in[1]
port 182 nsew signal input
flabel metal2 s 196778 -960 196890 480 0 FreeSans 448 90 0 0 la_data_in[20]
port 183 nsew signal input
flabel metal2 s 200274 -960 200386 480 0 FreeSans 448 90 0 0 la_data_in[21]
port 184 nsew signal input
flabel metal2 s 203862 -960 203974 480 0 FreeSans 448 90 0 0 la_data_in[22]
port 185 nsew signal input
flabel metal2 s 207358 -960 207470 480 0 FreeSans 448 90 0 0 la_data_in[23]
port 186 nsew signal input
flabel metal2 s 210946 -960 211058 480 0 FreeSans 448 90 0 0 la_data_in[24]
port 187 nsew signal input
flabel metal2 s 214442 -960 214554 480 0 FreeSans 448 90 0 0 la_data_in[25]
port 188 nsew signal input
flabel metal2 s 218030 -960 218142 480 0 FreeSans 448 90 0 0 la_data_in[26]
port 189 nsew signal input
flabel metal2 s 221526 -960 221638 480 0 FreeSans 448 90 0 0 la_data_in[27]
port 190 nsew signal input
flabel metal2 s 225114 -960 225226 480 0 FreeSans 448 90 0 0 la_data_in[28]
port 191 nsew signal input
flabel metal2 s 228702 -960 228814 480 0 FreeSans 448 90 0 0 la_data_in[29]
port 192 nsew signal input
flabel metal2 s 132930 -960 133042 480 0 FreeSans 448 90 0 0 la_data_in[2]
port 193 nsew signal input
flabel metal2 s 232198 -960 232310 480 0 FreeSans 448 90 0 0 la_data_in[30]
port 194 nsew signal input
flabel metal2 s 235786 -960 235898 480 0 FreeSans 448 90 0 0 la_data_in[31]
port 195 nsew signal input
flabel metal2 s 239282 -960 239394 480 0 FreeSans 448 90 0 0 la_data_in[32]
port 196 nsew signal input
flabel metal2 s 242870 -960 242982 480 0 FreeSans 448 90 0 0 la_data_in[33]
port 197 nsew signal input
flabel metal2 s 246366 -960 246478 480 0 FreeSans 448 90 0 0 la_data_in[34]
port 198 nsew signal input
flabel metal2 s 249954 -960 250066 480 0 FreeSans 448 90 0 0 la_data_in[35]
port 199 nsew signal input
flabel metal2 s 253450 -960 253562 480 0 FreeSans 448 90 0 0 la_data_in[36]
port 200 nsew signal input
flabel metal2 s 257038 -960 257150 480 0 FreeSans 448 90 0 0 la_data_in[37]
port 201 nsew signal input
flabel metal2 s 260626 -960 260738 480 0 FreeSans 448 90 0 0 la_data_in[38]
port 202 nsew signal input
flabel metal2 s 264122 -960 264234 480 0 FreeSans 448 90 0 0 la_data_in[39]
port 203 nsew signal input
flabel metal2 s 136426 -960 136538 480 0 FreeSans 448 90 0 0 la_data_in[3]
port 204 nsew signal input
flabel metal2 s 267710 -960 267822 480 0 FreeSans 448 90 0 0 la_data_in[40]
port 205 nsew signal input
flabel metal2 s 271206 -960 271318 480 0 FreeSans 448 90 0 0 la_data_in[41]
port 206 nsew signal input
flabel metal2 s 274794 -960 274906 480 0 FreeSans 448 90 0 0 la_data_in[42]
port 207 nsew signal input
flabel metal2 s 278290 -960 278402 480 0 FreeSans 448 90 0 0 la_data_in[43]
port 208 nsew signal input
flabel metal2 s 281878 -960 281990 480 0 FreeSans 448 90 0 0 la_data_in[44]
port 209 nsew signal input
flabel metal2 s 285374 -960 285486 480 0 FreeSans 448 90 0 0 la_data_in[45]
port 210 nsew signal input
flabel metal2 s 288962 -960 289074 480 0 FreeSans 448 90 0 0 la_data_in[46]
port 211 nsew signal input
flabel metal2 s 292550 -960 292662 480 0 FreeSans 448 90 0 0 la_data_in[47]
port 212 nsew signal input
flabel metal2 s 296046 -960 296158 480 0 FreeSans 448 90 0 0 la_data_in[48]
port 213 nsew signal input
flabel metal2 s 299634 -960 299746 480 0 FreeSans 448 90 0 0 la_data_in[49]
port 214 nsew signal input
flabel metal2 s 140014 -960 140126 480 0 FreeSans 448 90 0 0 la_data_in[4]
port 215 nsew signal input
flabel metal2 s 303130 -960 303242 480 0 FreeSans 448 90 0 0 la_data_in[50]
port 216 nsew signal input
flabel metal2 s 306718 -960 306830 480 0 FreeSans 448 90 0 0 la_data_in[51]
port 217 nsew signal input
flabel metal2 s 310214 -960 310326 480 0 FreeSans 448 90 0 0 la_data_in[52]
port 218 nsew signal input
flabel metal2 s 313802 -960 313914 480 0 FreeSans 448 90 0 0 la_data_in[53]
port 219 nsew signal input
flabel metal2 s 317298 -960 317410 480 0 FreeSans 448 90 0 0 la_data_in[54]
port 220 nsew signal input
flabel metal2 s 320886 -960 320998 480 0 FreeSans 448 90 0 0 la_data_in[55]
port 221 nsew signal input
flabel metal2 s 324382 -960 324494 480 0 FreeSans 448 90 0 0 la_data_in[56]
port 222 nsew signal input
flabel metal2 s 327970 -960 328082 480 0 FreeSans 448 90 0 0 la_data_in[57]
port 223 nsew signal input
flabel metal2 s 331558 -960 331670 480 0 FreeSans 448 90 0 0 la_data_in[58]
port 224 nsew signal input
flabel metal2 s 335054 -960 335166 480 0 FreeSans 448 90 0 0 la_data_in[59]
port 225 nsew signal input
flabel metal2 s 143510 -960 143622 480 0 FreeSans 448 90 0 0 la_data_in[5]
port 226 nsew signal input
flabel metal2 s 338642 -960 338754 480 0 FreeSans 448 90 0 0 la_data_in[60]
port 227 nsew signal input
flabel metal2 s 342138 -960 342250 480 0 FreeSans 448 90 0 0 la_data_in[61]
port 228 nsew signal input
flabel metal2 s 345726 -960 345838 480 0 FreeSans 448 90 0 0 la_data_in[62]
port 229 nsew signal input
flabel metal2 s 349222 -960 349334 480 0 FreeSans 448 90 0 0 la_data_in[63]
port 230 nsew signal input
flabel metal2 s 352810 -960 352922 480 0 FreeSans 448 90 0 0 la_data_in[64]
port 231 nsew signal input
flabel metal2 s 356306 -960 356418 480 0 FreeSans 448 90 0 0 la_data_in[65]
port 232 nsew signal input
flabel metal2 s 359894 -960 360006 480 0 FreeSans 448 90 0 0 la_data_in[66]
port 233 nsew signal input
flabel metal2 s 363482 -960 363594 480 0 FreeSans 448 90 0 0 la_data_in[67]
port 234 nsew signal input
flabel metal2 s 366978 -960 367090 480 0 FreeSans 448 90 0 0 la_data_in[68]
port 235 nsew signal input
flabel metal2 s 370566 -960 370678 480 0 FreeSans 448 90 0 0 la_data_in[69]
port 236 nsew signal input
flabel metal2 s 147098 -960 147210 480 0 FreeSans 448 90 0 0 la_data_in[6]
port 237 nsew signal input
flabel metal2 s 374062 -960 374174 480 0 FreeSans 448 90 0 0 la_data_in[70]
port 238 nsew signal input
flabel metal2 s 377650 -960 377762 480 0 FreeSans 448 90 0 0 la_data_in[71]
port 239 nsew signal input
flabel metal2 s 381146 -960 381258 480 0 FreeSans 448 90 0 0 la_data_in[72]
port 240 nsew signal input
flabel metal2 s 384734 -960 384846 480 0 FreeSans 448 90 0 0 la_data_in[73]
port 241 nsew signal input
flabel metal2 s 388230 -960 388342 480 0 FreeSans 448 90 0 0 la_data_in[74]
port 242 nsew signal input
flabel metal2 s 391818 -960 391930 480 0 FreeSans 448 90 0 0 la_data_in[75]
port 243 nsew signal input
flabel metal2 s 395314 -960 395426 480 0 FreeSans 448 90 0 0 la_data_in[76]
port 244 nsew signal input
flabel metal2 s 398902 -960 399014 480 0 FreeSans 448 90 0 0 la_data_in[77]
port 245 nsew signal input
flabel metal2 s 402490 -960 402602 480 0 FreeSans 448 90 0 0 la_data_in[78]
port 246 nsew signal input
flabel metal2 s 405986 -960 406098 480 0 FreeSans 448 90 0 0 la_data_in[79]
port 247 nsew signal input
flabel metal2 s 150594 -960 150706 480 0 FreeSans 448 90 0 0 la_data_in[7]
port 248 nsew signal input
flabel metal2 s 409574 -960 409686 480 0 FreeSans 448 90 0 0 la_data_in[80]
port 249 nsew signal input
flabel metal2 s 413070 -960 413182 480 0 FreeSans 448 90 0 0 la_data_in[81]
port 250 nsew signal input
flabel metal2 s 416658 -960 416770 480 0 FreeSans 448 90 0 0 la_data_in[82]
port 251 nsew signal input
flabel metal2 s 420154 -960 420266 480 0 FreeSans 448 90 0 0 la_data_in[83]
port 252 nsew signal input
flabel metal2 s 423742 -960 423854 480 0 FreeSans 448 90 0 0 la_data_in[84]
port 253 nsew signal input
flabel metal2 s 427238 -960 427350 480 0 FreeSans 448 90 0 0 la_data_in[85]
port 254 nsew signal input
flabel metal2 s 430826 -960 430938 480 0 FreeSans 448 90 0 0 la_data_in[86]
port 255 nsew signal input
flabel metal2 s 434414 -960 434526 480 0 FreeSans 448 90 0 0 la_data_in[87]
port 256 nsew signal input
flabel metal2 s 437910 -960 438022 480 0 FreeSans 448 90 0 0 la_data_in[88]
port 257 nsew signal input
flabel metal2 s 441498 -960 441610 480 0 FreeSans 448 90 0 0 la_data_in[89]
port 258 nsew signal input
flabel metal2 s 154182 -960 154294 480 0 FreeSans 448 90 0 0 la_data_in[8]
port 259 nsew signal input
flabel metal2 s 444994 -960 445106 480 0 FreeSans 448 90 0 0 la_data_in[90]
port 260 nsew signal input
flabel metal2 s 448582 -960 448694 480 0 FreeSans 448 90 0 0 la_data_in[91]
port 261 nsew signal input
flabel metal2 s 452078 -960 452190 480 0 FreeSans 448 90 0 0 la_data_in[92]
port 262 nsew signal input
flabel metal2 s 455666 -960 455778 480 0 FreeSans 448 90 0 0 la_data_in[93]
port 263 nsew signal input
flabel metal2 s 459162 -960 459274 480 0 FreeSans 448 90 0 0 la_data_in[94]
port 264 nsew signal input
flabel metal2 s 462750 -960 462862 480 0 FreeSans 448 90 0 0 la_data_in[95]
port 265 nsew signal input
flabel metal2 s 466246 -960 466358 480 0 FreeSans 448 90 0 0 la_data_in[96]
port 266 nsew signal input
flabel metal2 s 469834 -960 469946 480 0 FreeSans 448 90 0 0 la_data_in[97]
port 267 nsew signal input
flabel metal2 s 473422 -960 473534 480 0 FreeSans 448 90 0 0 la_data_in[98]
port 268 nsew signal input
flabel metal2 s 476918 -960 477030 480 0 FreeSans 448 90 0 0 la_data_in[99]
port 269 nsew signal input
flabel metal2 s 157770 -960 157882 480 0 FreeSans 448 90 0 0 la_data_in[9]
port 270 nsew signal input
flabel metal2 s 126950 -960 127062 480 0 FreeSans 448 90 0 0 la_data_out[0]
port 271 nsew signal tristate
flabel metal2 s 481702 -960 481814 480 0 FreeSans 448 90 0 0 la_data_out[100]
port 272 nsew signal tristate
flabel metal2 s 485198 -960 485310 480 0 FreeSans 448 90 0 0 la_data_out[101]
port 273 nsew signal tristate
flabel metal2 s 488786 -960 488898 480 0 FreeSans 448 90 0 0 la_data_out[102]
port 274 nsew signal tristate
flabel metal2 s 492282 -960 492394 480 0 FreeSans 448 90 0 0 la_data_out[103]
port 275 nsew signal tristate
flabel metal2 s 495870 -960 495982 480 0 FreeSans 448 90 0 0 la_data_out[104]
port 276 nsew signal tristate
flabel metal2 s 499366 -960 499478 480 0 FreeSans 448 90 0 0 la_data_out[105]
port 277 nsew signal tristate
flabel metal2 s 502954 -960 503066 480 0 FreeSans 448 90 0 0 la_data_out[106]
port 278 nsew signal tristate
flabel metal2 s 506450 -960 506562 480 0 FreeSans 448 90 0 0 la_data_out[107]
port 279 nsew signal tristate
flabel metal2 s 510038 -960 510150 480 0 FreeSans 448 90 0 0 la_data_out[108]
port 280 nsew signal tristate
flabel metal2 s 513534 -960 513646 480 0 FreeSans 448 90 0 0 la_data_out[109]
port 281 nsew signal tristate
flabel metal2 s 162462 -960 162574 480 0 FreeSans 448 90 0 0 la_data_out[10]
port 282 nsew signal tristate
flabel metal2 s 517122 -960 517234 480 0 FreeSans 448 90 0 0 la_data_out[110]
port 283 nsew signal tristate
flabel metal2 s 520710 -960 520822 480 0 FreeSans 448 90 0 0 la_data_out[111]
port 284 nsew signal tristate
flabel metal2 s 524206 -960 524318 480 0 FreeSans 448 90 0 0 la_data_out[112]
port 285 nsew signal tristate
flabel metal2 s 527794 -960 527906 480 0 FreeSans 448 90 0 0 la_data_out[113]
port 286 nsew signal tristate
flabel metal2 s 531290 -960 531402 480 0 FreeSans 448 90 0 0 la_data_out[114]
port 287 nsew signal tristate
flabel metal2 s 534878 -960 534990 480 0 FreeSans 448 90 0 0 la_data_out[115]
port 288 nsew signal tristate
flabel metal2 s 538374 -960 538486 480 0 FreeSans 448 90 0 0 la_data_out[116]
port 289 nsew signal tristate
flabel metal2 s 541962 -960 542074 480 0 FreeSans 448 90 0 0 la_data_out[117]
port 290 nsew signal tristate
flabel metal2 s 545458 -960 545570 480 0 FreeSans 448 90 0 0 la_data_out[118]
port 291 nsew signal tristate
flabel metal2 s 549046 -960 549158 480 0 FreeSans 448 90 0 0 la_data_out[119]
port 292 nsew signal tristate
flabel metal2 s 166050 -960 166162 480 0 FreeSans 448 90 0 0 la_data_out[11]
port 293 nsew signal tristate
flabel metal2 s 552634 -960 552746 480 0 FreeSans 448 90 0 0 la_data_out[120]
port 294 nsew signal tristate
flabel metal2 s 556130 -960 556242 480 0 FreeSans 448 90 0 0 la_data_out[121]
port 295 nsew signal tristate
flabel metal2 s 559718 -960 559830 480 0 FreeSans 448 90 0 0 la_data_out[122]
port 296 nsew signal tristate
flabel metal2 s 563214 -960 563326 480 0 FreeSans 448 90 0 0 la_data_out[123]
port 297 nsew signal tristate
flabel metal2 s 566802 -960 566914 480 0 FreeSans 448 90 0 0 la_data_out[124]
port 298 nsew signal tristate
flabel metal2 s 570298 -960 570410 480 0 FreeSans 448 90 0 0 la_data_out[125]
port 299 nsew signal tristate
flabel metal2 s 573886 -960 573998 480 0 FreeSans 448 90 0 0 la_data_out[126]
port 300 nsew signal tristate
flabel metal2 s 577382 -960 577494 480 0 FreeSans 448 90 0 0 la_data_out[127]
port 301 nsew signal tristate
flabel metal2 s 169546 -960 169658 480 0 FreeSans 448 90 0 0 la_data_out[12]
port 302 nsew signal tristate
flabel metal2 s 173134 -960 173246 480 0 FreeSans 448 90 0 0 la_data_out[13]
port 303 nsew signal tristate
flabel metal2 s 176630 -960 176742 480 0 FreeSans 448 90 0 0 la_data_out[14]
port 304 nsew signal tristate
flabel metal2 s 180218 -960 180330 480 0 FreeSans 448 90 0 0 la_data_out[15]
port 305 nsew signal tristate
flabel metal2 s 183714 -960 183826 480 0 FreeSans 448 90 0 0 la_data_out[16]
port 306 nsew signal tristate
flabel metal2 s 187302 -960 187414 480 0 FreeSans 448 90 0 0 la_data_out[17]
port 307 nsew signal tristate
flabel metal2 s 190798 -960 190910 480 0 FreeSans 448 90 0 0 la_data_out[18]
port 308 nsew signal tristate
flabel metal2 s 194386 -960 194498 480 0 FreeSans 448 90 0 0 la_data_out[19]
port 309 nsew signal tristate
flabel metal2 s 130538 -960 130650 480 0 FreeSans 448 90 0 0 la_data_out[1]
port 310 nsew signal tristate
flabel metal2 s 197882 -960 197994 480 0 FreeSans 448 90 0 0 la_data_out[20]
port 311 nsew signal tristate
flabel metal2 s 201470 -960 201582 480 0 FreeSans 448 90 0 0 la_data_out[21]
port 312 nsew signal tristate
flabel metal2 s 205058 -960 205170 480 0 FreeSans 448 90 0 0 la_data_out[22]
port 313 nsew signal tristate
flabel metal2 s 208554 -960 208666 480 0 FreeSans 448 90 0 0 la_data_out[23]
port 314 nsew signal tristate
flabel metal2 s 212142 -960 212254 480 0 FreeSans 448 90 0 0 la_data_out[24]
port 315 nsew signal tristate
flabel metal2 s 215638 -960 215750 480 0 FreeSans 448 90 0 0 la_data_out[25]
port 316 nsew signal tristate
flabel metal2 s 219226 -960 219338 480 0 FreeSans 448 90 0 0 la_data_out[26]
port 317 nsew signal tristate
flabel metal2 s 222722 -960 222834 480 0 FreeSans 448 90 0 0 la_data_out[27]
port 318 nsew signal tristate
flabel metal2 s 226310 -960 226422 480 0 FreeSans 448 90 0 0 la_data_out[28]
port 319 nsew signal tristate
flabel metal2 s 229806 -960 229918 480 0 FreeSans 448 90 0 0 la_data_out[29]
port 320 nsew signal tristate
flabel metal2 s 134126 -960 134238 480 0 FreeSans 448 90 0 0 la_data_out[2]
port 321 nsew signal tristate
flabel metal2 s 233394 -960 233506 480 0 FreeSans 448 90 0 0 la_data_out[30]
port 322 nsew signal tristate
flabel metal2 s 236982 -960 237094 480 0 FreeSans 448 90 0 0 la_data_out[31]
port 323 nsew signal tristate
flabel metal2 s 240478 -960 240590 480 0 FreeSans 448 90 0 0 la_data_out[32]
port 324 nsew signal tristate
flabel metal2 s 244066 -960 244178 480 0 FreeSans 448 90 0 0 la_data_out[33]
port 325 nsew signal tristate
flabel metal2 s 247562 -960 247674 480 0 FreeSans 448 90 0 0 la_data_out[34]
port 326 nsew signal tristate
flabel metal2 s 251150 -960 251262 480 0 FreeSans 448 90 0 0 la_data_out[35]
port 327 nsew signal tristate
flabel metal2 s 254646 -960 254758 480 0 FreeSans 448 90 0 0 la_data_out[36]
port 328 nsew signal tristate
flabel metal2 s 258234 -960 258346 480 0 FreeSans 448 90 0 0 la_data_out[37]
port 329 nsew signal tristate
flabel metal2 s 261730 -960 261842 480 0 FreeSans 448 90 0 0 la_data_out[38]
port 330 nsew signal tristate
flabel metal2 s 265318 -960 265430 480 0 FreeSans 448 90 0 0 la_data_out[39]
port 331 nsew signal tristate
flabel metal2 s 137622 -960 137734 480 0 FreeSans 448 90 0 0 la_data_out[3]
port 332 nsew signal tristate
flabel metal2 s 268814 -960 268926 480 0 FreeSans 448 90 0 0 la_data_out[40]
port 333 nsew signal tristate
flabel metal2 s 272402 -960 272514 480 0 FreeSans 448 90 0 0 la_data_out[41]
port 334 nsew signal tristate
flabel metal2 s 275990 -960 276102 480 0 FreeSans 448 90 0 0 la_data_out[42]
port 335 nsew signal tristate
flabel metal2 s 279486 -960 279598 480 0 FreeSans 448 90 0 0 la_data_out[43]
port 336 nsew signal tristate
flabel metal2 s 283074 -960 283186 480 0 FreeSans 448 90 0 0 la_data_out[44]
port 337 nsew signal tristate
flabel metal2 s 286570 -960 286682 480 0 FreeSans 448 90 0 0 la_data_out[45]
port 338 nsew signal tristate
flabel metal2 s 290158 -960 290270 480 0 FreeSans 448 90 0 0 la_data_out[46]
port 339 nsew signal tristate
flabel metal2 s 293654 -960 293766 480 0 FreeSans 448 90 0 0 la_data_out[47]
port 340 nsew signal tristate
flabel metal2 s 297242 -960 297354 480 0 FreeSans 448 90 0 0 la_data_out[48]
port 341 nsew signal tristate
flabel metal2 s 300738 -960 300850 480 0 FreeSans 448 90 0 0 la_data_out[49]
port 342 nsew signal tristate
flabel metal2 s 141210 -960 141322 480 0 FreeSans 448 90 0 0 la_data_out[4]
port 343 nsew signal tristate
flabel metal2 s 304326 -960 304438 480 0 FreeSans 448 90 0 0 la_data_out[50]
port 344 nsew signal tristate
flabel metal2 s 307914 -960 308026 480 0 FreeSans 448 90 0 0 la_data_out[51]
port 345 nsew signal tristate
flabel metal2 s 311410 -960 311522 480 0 FreeSans 448 90 0 0 la_data_out[52]
port 346 nsew signal tristate
flabel metal2 s 314998 -960 315110 480 0 FreeSans 448 90 0 0 la_data_out[53]
port 347 nsew signal tristate
flabel metal2 s 318494 -960 318606 480 0 FreeSans 448 90 0 0 la_data_out[54]
port 348 nsew signal tristate
flabel metal2 s 322082 -960 322194 480 0 FreeSans 448 90 0 0 la_data_out[55]
port 349 nsew signal tristate
flabel metal2 s 325578 -960 325690 480 0 FreeSans 448 90 0 0 la_data_out[56]
port 350 nsew signal tristate
flabel metal2 s 329166 -960 329278 480 0 FreeSans 448 90 0 0 la_data_out[57]
port 351 nsew signal tristate
flabel metal2 s 332662 -960 332774 480 0 FreeSans 448 90 0 0 la_data_out[58]
port 352 nsew signal tristate
flabel metal2 s 336250 -960 336362 480 0 FreeSans 448 90 0 0 la_data_out[59]
port 353 nsew signal tristate
flabel metal2 s 144706 -960 144818 480 0 FreeSans 448 90 0 0 la_data_out[5]
port 354 nsew signal tristate
flabel metal2 s 339838 -960 339950 480 0 FreeSans 448 90 0 0 la_data_out[60]
port 355 nsew signal tristate
flabel metal2 s 343334 -960 343446 480 0 FreeSans 448 90 0 0 la_data_out[61]
port 356 nsew signal tristate
flabel metal2 s 346922 -960 347034 480 0 FreeSans 448 90 0 0 la_data_out[62]
port 357 nsew signal tristate
flabel metal2 s 350418 -960 350530 480 0 FreeSans 448 90 0 0 la_data_out[63]
port 358 nsew signal tristate
flabel metal2 s 354006 -960 354118 480 0 FreeSans 448 90 0 0 la_data_out[64]
port 359 nsew signal tristate
flabel metal2 s 357502 -960 357614 480 0 FreeSans 448 90 0 0 la_data_out[65]
port 360 nsew signal tristate
flabel metal2 s 361090 -960 361202 480 0 FreeSans 448 90 0 0 la_data_out[66]
port 361 nsew signal tristate
flabel metal2 s 364586 -960 364698 480 0 FreeSans 448 90 0 0 la_data_out[67]
port 362 nsew signal tristate
flabel metal2 s 368174 -960 368286 480 0 FreeSans 448 90 0 0 la_data_out[68]
port 363 nsew signal tristate
flabel metal2 s 371670 -960 371782 480 0 FreeSans 448 90 0 0 la_data_out[69]
port 364 nsew signal tristate
flabel metal2 s 148294 -960 148406 480 0 FreeSans 448 90 0 0 la_data_out[6]
port 365 nsew signal tristate
flabel metal2 s 375258 -960 375370 480 0 FreeSans 448 90 0 0 la_data_out[70]
port 366 nsew signal tristate
flabel metal2 s 378846 -960 378958 480 0 FreeSans 448 90 0 0 la_data_out[71]
port 367 nsew signal tristate
flabel metal2 s 382342 -960 382454 480 0 FreeSans 448 90 0 0 la_data_out[72]
port 368 nsew signal tristate
flabel metal2 s 385930 -960 386042 480 0 FreeSans 448 90 0 0 la_data_out[73]
port 369 nsew signal tristate
flabel metal2 s 389426 -960 389538 480 0 FreeSans 448 90 0 0 la_data_out[74]
port 370 nsew signal tristate
flabel metal2 s 393014 -960 393126 480 0 FreeSans 448 90 0 0 la_data_out[75]
port 371 nsew signal tristate
flabel metal2 s 396510 -960 396622 480 0 FreeSans 448 90 0 0 la_data_out[76]
port 372 nsew signal tristate
flabel metal2 s 400098 -960 400210 480 0 FreeSans 448 90 0 0 la_data_out[77]
port 373 nsew signal tristate
flabel metal2 s 403594 -960 403706 480 0 FreeSans 448 90 0 0 la_data_out[78]
port 374 nsew signal tristate
flabel metal2 s 407182 -960 407294 480 0 FreeSans 448 90 0 0 la_data_out[79]
port 375 nsew signal tristate
flabel metal2 s 151790 -960 151902 480 0 FreeSans 448 90 0 0 la_data_out[7]
port 376 nsew signal tristate
flabel metal2 s 410770 -960 410882 480 0 FreeSans 448 90 0 0 la_data_out[80]
port 377 nsew signal tristate
flabel metal2 s 414266 -960 414378 480 0 FreeSans 448 90 0 0 la_data_out[81]
port 378 nsew signal tristate
flabel metal2 s 417854 -960 417966 480 0 FreeSans 448 90 0 0 la_data_out[82]
port 379 nsew signal tristate
flabel metal2 s 421350 -960 421462 480 0 FreeSans 448 90 0 0 la_data_out[83]
port 380 nsew signal tristate
flabel metal2 s 424938 -960 425050 480 0 FreeSans 448 90 0 0 la_data_out[84]
port 381 nsew signal tristate
flabel metal2 s 428434 -960 428546 480 0 FreeSans 448 90 0 0 la_data_out[85]
port 382 nsew signal tristate
flabel metal2 s 432022 -960 432134 480 0 FreeSans 448 90 0 0 la_data_out[86]
port 383 nsew signal tristate
flabel metal2 s 435518 -960 435630 480 0 FreeSans 448 90 0 0 la_data_out[87]
port 384 nsew signal tristate
flabel metal2 s 439106 -960 439218 480 0 FreeSans 448 90 0 0 la_data_out[88]
port 385 nsew signal tristate
flabel metal2 s 442602 -960 442714 480 0 FreeSans 448 90 0 0 la_data_out[89]
port 386 nsew signal tristate
flabel metal2 s 155378 -960 155490 480 0 FreeSans 448 90 0 0 la_data_out[8]
port 387 nsew signal tristate
flabel metal2 s 446190 -960 446302 480 0 FreeSans 448 90 0 0 la_data_out[90]
port 388 nsew signal tristate
flabel metal2 s 449778 -960 449890 480 0 FreeSans 448 90 0 0 la_data_out[91]
port 389 nsew signal tristate
flabel metal2 s 453274 -960 453386 480 0 FreeSans 448 90 0 0 la_data_out[92]
port 390 nsew signal tristate
flabel metal2 s 456862 -960 456974 480 0 FreeSans 448 90 0 0 la_data_out[93]
port 391 nsew signal tristate
flabel metal2 s 460358 -960 460470 480 0 FreeSans 448 90 0 0 la_data_out[94]
port 392 nsew signal tristate
flabel metal2 s 463946 -960 464058 480 0 FreeSans 448 90 0 0 la_data_out[95]
port 393 nsew signal tristate
flabel metal2 s 467442 -960 467554 480 0 FreeSans 448 90 0 0 la_data_out[96]
port 394 nsew signal tristate
flabel metal2 s 471030 -960 471142 480 0 FreeSans 448 90 0 0 la_data_out[97]
port 395 nsew signal tristate
flabel metal2 s 474526 -960 474638 480 0 FreeSans 448 90 0 0 la_data_out[98]
port 396 nsew signal tristate
flabel metal2 s 478114 -960 478226 480 0 FreeSans 448 90 0 0 la_data_out[99]
port 397 nsew signal tristate
flabel metal2 s 158874 -960 158986 480 0 FreeSans 448 90 0 0 la_data_out[9]
port 398 nsew signal tristate
flabel metal2 s 128146 -960 128258 480 0 FreeSans 448 90 0 0 la_oenb[0]
port 399 nsew signal input
flabel metal2 s 482806 -960 482918 480 0 FreeSans 448 90 0 0 la_oenb[100]
port 400 nsew signal input
flabel metal2 s 486394 -960 486506 480 0 FreeSans 448 90 0 0 la_oenb[101]
port 401 nsew signal input
flabel metal2 s 489890 -960 490002 480 0 FreeSans 448 90 0 0 la_oenb[102]
port 402 nsew signal input
flabel metal2 s 493478 -960 493590 480 0 FreeSans 448 90 0 0 la_oenb[103]
port 403 nsew signal input
flabel metal2 s 497066 -960 497178 480 0 FreeSans 448 90 0 0 la_oenb[104]
port 404 nsew signal input
flabel metal2 s 500562 -960 500674 480 0 FreeSans 448 90 0 0 la_oenb[105]
port 405 nsew signal input
flabel metal2 s 504150 -960 504262 480 0 FreeSans 448 90 0 0 la_oenb[106]
port 406 nsew signal input
flabel metal2 s 507646 -960 507758 480 0 FreeSans 448 90 0 0 la_oenb[107]
port 407 nsew signal input
flabel metal2 s 511234 -960 511346 480 0 FreeSans 448 90 0 0 la_oenb[108]
port 408 nsew signal input
flabel metal2 s 514730 -960 514842 480 0 FreeSans 448 90 0 0 la_oenb[109]
port 409 nsew signal input
flabel metal2 s 163658 -960 163770 480 0 FreeSans 448 90 0 0 la_oenb[10]
port 410 nsew signal input
flabel metal2 s 518318 -960 518430 480 0 FreeSans 448 90 0 0 la_oenb[110]
port 411 nsew signal input
flabel metal2 s 521814 -960 521926 480 0 FreeSans 448 90 0 0 la_oenb[111]
port 412 nsew signal input
flabel metal2 s 525402 -960 525514 480 0 FreeSans 448 90 0 0 la_oenb[112]
port 413 nsew signal input
flabel metal2 s 528990 -960 529102 480 0 FreeSans 448 90 0 0 la_oenb[113]
port 414 nsew signal input
flabel metal2 s 532486 -960 532598 480 0 FreeSans 448 90 0 0 la_oenb[114]
port 415 nsew signal input
flabel metal2 s 536074 -960 536186 480 0 FreeSans 448 90 0 0 la_oenb[115]
port 416 nsew signal input
flabel metal2 s 539570 -960 539682 480 0 FreeSans 448 90 0 0 la_oenb[116]
port 417 nsew signal input
flabel metal2 s 543158 -960 543270 480 0 FreeSans 448 90 0 0 la_oenb[117]
port 418 nsew signal input
flabel metal2 s 546654 -960 546766 480 0 FreeSans 448 90 0 0 la_oenb[118]
port 419 nsew signal input
flabel metal2 s 550242 -960 550354 480 0 FreeSans 448 90 0 0 la_oenb[119]
port 420 nsew signal input
flabel metal2 s 167154 -960 167266 480 0 FreeSans 448 90 0 0 la_oenb[11]
port 421 nsew signal input
flabel metal2 s 553738 -960 553850 480 0 FreeSans 448 90 0 0 la_oenb[120]
port 422 nsew signal input
flabel metal2 s 557326 -960 557438 480 0 FreeSans 448 90 0 0 la_oenb[121]
port 423 nsew signal input
flabel metal2 s 560822 -960 560934 480 0 FreeSans 448 90 0 0 la_oenb[122]
port 424 nsew signal input
flabel metal2 s 564410 -960 564522 480 0 FreeSans 448 90 0 0 la_oenb[123]
port 425 nsew signal input
flabel metal2 s 567998 -960 568110 480 0 FreeSans 448 90 0 0 la_oenb[124]
port 426 nsew signal input
flabel metal2 s 571494 -960 571606 480 0 FreeSans 448 90 0 0 la_oenb[125]
port 427 nsew signal input
flabel metal2 s 575082 -960 575194 480 0 FreeSans 448 90 0 0 la_oenb[126]
port 428 nsew signal input
flabel metal2 s 578578 -960 578690 480 0 FreeSans 448 90 0 0 la_oenb[127]
port 429 nsew signal input
flabel metal2 s 170742 -960 170854 480 0 FreeSans 448 90 0 0 la_oenb[12]
port 430 nsew signal input
flabel metal2 s 174238 -960 174350 480 0 FreeSans 448 90 0 0 la_oenb[13]
port 431 nsew signal input
flabel metal2 s 177826 -960 177938 480 0 FreeSans 448 90 0 0 la_oenb[14]
port 432 nsew signal input
flabel metal2 s 181414 -960 181526 480 0 FreeSans 448 90 0 0 la_oenb[15]
port 433 nsew signal input
flabel metal2 s 184910 -960 185022 480 0 FreeSans 448 90 0 0 la_oenb[16]
port 434 nsew signal input
flabel metal2 s 188498 -960 188610 480 0 FreeSans 448 90 0 0 la_oenb[17]
port 435 nsew signal input
flabel metal2 s 191994 -960 192106 480 0 FreeSans 448 90 0 0 la_oenb[18]
port 436 nsew signal input
flabel metal2 s 195582 -960 195694 480 0 FreeSans 448 90 0 0 la_oenb[19]
port 437 nsew signal input
flabel metal2 s 131734 -960 131846 480 0 FreeSans 448 90 0 0 la_oenb[1]
port 438 nsew signal input
flabel metal2 s 199078 -960 199190 480 0 FreeSans 448 90 0 0 la_oenb[20]
port 439 nsew signal input
flabel metal2 s 202666 -960 202778 480 0 FreeSans 448 90 0 0 la_oenb[21]
port 440 nsew signal input
flabel metal2 s 206162 -960 206274 480 0 FreeSans 448 90 0 0 la_oenb[22]
port 441 nsew signal input
flabel metal2 s 209750 -960 209862 480 0 FreeSans 448 90 0 0 la_oenb[23]
port 442 nsew signal input
flabel metal2 s 213338 -960 213450 480 0 FreeSans 448 90 0 0 la_oenb[24]
port 443 nsew signal input
flabel metal2 s 216834 -960 216946 480 0 FreeSans 448 90 0 0 la_oenb[25]
port 444 nsew signal input
flabel metal2 s 220422 -960 220534 480 0 FreeSans 448 90 0 0 la_oenb[26]
port 445 nsew signal input
flabel metal2 s 223918 -960 224030 480 0 FreeSans 448 90 0 0 la_oenb[27]
port 446 nsew signal input
flabel metal2 s 227506 -960 227618 480 0 FreeSans 448 90 0 0 la_oenb[28]
port 447 nsew signal input
flabel metal2 s 231002 -960 231114 480 0 FreeSans 448 90 0 0 la_oenb[29]
port 448 nsew signal input
flabel metal2 s 135230 -960 135342 480 0 FreeSans 448 90 0 0 la_oenb[2]
port 449 nsew signal input
flabel metal2 s 234590 -960 234702 480 0 FreeSans 448 90 0 0 la_oenb[30]
port 450 nsew signal input
flabel metal2 s 238086 -960 238198 480 0 FreeSans 448 90 0 0 la_oenb[31]
port 451 nsew signal input
flabel metal2 s 241674 -960 241786 480 0 FreeSans 448 90 0 0 la_oenb[32]
port 452 nsew signal input
flabel metal2 s 245170 -960 245282 480 0 FreeSans 448 90 0 0 la_oenb[33]
port 453 nsew signal input
flabel metal2 s 248758 -960 248870 480 0 FreeSans 448 90 0 0 la_oenb[34]
port 454 nsew signal input
flabel metal2 s 252346 -960 252458 480 0 FreeSans 448 90 0 0 la_oenb[35]
port 455 nsew signal input
flabel metal2 s 255842 -960 255954 480 0 FreeSans 448 90 0 0 la_oenb[36]
port 456 nsew signal input
flabel metal2 s 259430 -960 259542 480 0 FreeSans 448 90 0 0 la_oenb[37]
port 457 nsew signal input
flabel metal2 s 262926 -960 263038 480 0 FreeSans 448 90 0 0 la_oenb[38]
port 458 nsew signal input
flabel metal2 s 266514 -960 266626 480 0 FreeSans 448 90 0 0 la_oenb[39]
port 459 nsew signal input
flabel metal2 s 138818 -960 138930 480 0 FreeSans 448 90 0 0 la_oenb[3]
port 460 nsew signal input
flabel metal2 s 270010 -960 270122 480 0 FreeSans 448 90 0 0 la_oenb[40]
port 461 nsew signal input
flabel metal2 s 273598 -960 273710 480 0 FreeSans 448 90 0 0 la_oenb[41]
port 462 nsew signal input
flabel metal2 s 277094 -960 277206 480 0 FreeSans 448 90 0 0 la_oenb[42]
port 463 nsew signal input
flabel metal2 s 280682 -960 280794 480 0 FreeSans 448 90 0 0 la_oenb[43]
port 464 nsew signal input
flabel metal2 s 284270 -960 284382 480 0 FreeSans 448 90 0 0 la_oenb[44]
port 465 nsew signal input
flabel metal2 s 287766 -960 287878 480 0 FreeSans 448 90 0 0 la_oenb[45]
port 466 nsew signal input
flabel metal2 s 291354 -960 291466 480 0 FreeSans 448 90 0 0 la_oenb[46]
port 467 nsew signal input
flabel metal2 s 294850 -960 294962 480 0 FreeSans 448 90 0 0 la_oenb[47]
port 468 nsew signal input
flabel metal2 s 298438 -960 298550 480 0 FreeSans 448 90 0 0 la_oenb[48]
port 469 nsew signal input
flabel metal2 s 301934 -960 302046 480 0 FreeSans 448 90 0 0 la_oenb[49]
port 470 nsew signal input
flabel metal2 s 142406 -960 142518 480 0 FreeSans 448 90 0 0 la_oenb[4]
port 471 nsew signal input
flabel metal2 s 305522 -960 305634 480 0 FreeSans 448 90 0 0 la_oenb[50]
port 472 nsew signal input
flabel metal2 s 309018 -960 309130 480 0 FreeSans 448 90 0 0 la_oenb[51]
port 473 nsew signal input
flabel metal2 s 312606 -960 312718 480 0 FreeSans 448 90 0 0 la_oenb[52]
port 474 nsew signal input
flabel metal2 s 316194 -960 316306 480 0 FreeSans 448 90 0 0 la_oenb[53]
port 475 nsew signal input
flabel metal2 s 319690 -960 319802 480 0 FreeSans 448 90 0 0 la_oenb[54]
port 476 nsew signal input
flabel metal2 s 323278 -960 323390 480 0 FreeSans 448 90 0 0 la_oenb[55]
port 477 nsew signal input
flabel metal2 s 326774 -960 326886 480 0 FreeSans 448 90 0 0 la_oenb[56]
port 478 nsew signal input
flabel metal2 s 330362 -960 330474 480 0 FreeSans 448 90 0 0 la_oenb[57]
port 479 nsew signal input
flabel metal2 s 333858 -960 333970 480 0 FreeSans 448 90 0 0 la_oenb[58]
port 480 nsew signal input
flabel metal2 s 337446 -960 337558 480 0 FreeSans 448 90 0 0 la_oenb[59]
port 481 nsew signal input
flabel metal2 s 145902 -960 146014 480 0 FreeSans 448 90 0 0 la_oenb[5]
port 482 nsew signal input
flabel metal2 s 340942 -960 341054 480 0 FreeSans 448 90 0 0 la_oenb[60]
port 483 nsew signal input
flabel metal2 s 344530 -960 344642 480 0 FreeSans 448 90 0 0 la_oenb[61]
port 484 nsew signal input
flabel metal2 s 348026 -960 348138 480 0 FreeSans 448 90 0 0 la_oenb[62]
port 485 nsew signal input
flabel metal2 s 351614 -960 351726 480 0 FreeSans 448 90 0 0 la_oenb[63]
port 486 nsew signal input
flabel metal2 s 355202 -960 355314 480 0 FreeSans 448 90 0 0 la_oenb[64]
port 487 nsew signal input
flabel metal2 s 358698 -960 358810 480 0 FreeSans 448 90 0 0 la_oenb[65]
port 488 nsew signal input
flabel metal2 s 362286 -960 362398 480 0 FreeSans 448 90 0 0 la_oenb[66]
port 489 nsew signal input
flabel metal2 s 365782 -960 365894 480 0 FreeSans 448 90 0 0 la_oenb[67]
port 490 nsew signal input
flabel metal2 s 369370 -960 369482 480 0 FreeSans 448 90 0 0 la_oenb[68]
port 491 nsew signal input
flabel metal2 s 372866 -960 372978 480 0 FreeSans 448 90 0 0 la_oenb[69]
port 492 nsew signal input
flabel metal2 s 149490 -960 149602 480 0 FreeSans 448 90 0 0 la_oenb[6]
port 493 nsew signal input
flabel metal2 s 376454 -960 376566 480 0 FreeSans 448 90 0 0 la_oenb[70]
port 494 nsew signal input
flabel metal2 s 379950 -960 380062 480 0 FreeSans 448 90 0 0 la_oenb[71]
port 495 nsew signal input
flabel metal2 s 383538 -960 383650 480 0 FreeSans 448 90 0 0 la_oenb[72]
port 496 nsew signal input
flabel metal2 s 387126 -960 387238 480 0 FreeSans 448 90 0 0 la_oenb[73]
port 497 nsew signal input
flabel metal2 s 390622 -960 390734 480 0 FreeSans 448 90 0 0 la_oenb[74]
port 498 nsew signal input
flabel metal2 s 394210 -960 394322 480 0 FreeSans 448 90 0 0 la_oenb[75]
port 499 nsew signal input
flabel metal2 s 397706 -960 397818 480 0 FreeSans 448 90 0 0 la_oenb[76]
port 500 nsew signal input
flabel metal2 s 401294 -960 401406 480 0 FreeSans 448 90 0 0 la_oenb[77]
port 501 nsew signal input
flabel metal2 s 404790 -960 404902 480 0 FreeSans 448 90 0 0 la_oenb[78]
port 502 nsew signal input
flabel metal2 s 408378 -960 408490 480 0 FreeSans 448 90 0 0 la_oenb[79]
port 503 nsew signal input
flabel metal2 s 152986 -960 153098 480 0 FreeSans 448 90 0 0 la_oenb[7]
port 504 nsew signal input
flabel metal2 s 411874 -960 411986 480 0 FreeSans 448 90 0 0 la_oenb[80]
port 505 nsew signal input
flabel metal2 s 415462 -960 415574 480 0 FreeSans 448 90 0 0 la_oenb[81]
port 506 nsew signal input
flabel metal2 s 418958 -960 419070 480 0 FreeSans 448 90 0 0 la_oenb[82]
port 507 nsew signal input
flabel metal2 s 422546 -960 422658 480 0 FreeSans 448 90 0 0 la_oenb[83]
port 508 nsew signal input
flabel metal2 s 426134 -960 426246 480 0 FreeSans 448 90 0 0 la_oenb[84]
port 509 nsew signal input
flabel metal2 s 429630 -960 429742 480 0 FreeSans 448 90 0 0 la_oenb[85]
port 510 nsew signal input
flabel metal2 s 433218 -960 433330 480 0 FreeSans 448 90 0 0 la_oenb[86]
port 511 nsew signal input
flabel metal2 s 436714 -960 436826 480 0 FreeSans 448 90 0 0 la_oenb[87]
port 512 nsew signal input
flabel metal2 s 440302 -960 440414 480 0 FreeSans 448 90 0 0 la_oenb[88]
port 513 nsew signal input
flabel metal2 s 443798 -960 443910 480 0 FreeSans 448 90 0 0 la_oenb[89]
port 514 nsew signal input
flabel metal2 s 156574 -960 156686 480 0 FreeSans 448 90 0 0 la_oenb[8]
port 515 nsew signal input
flabel metal2 s 447386 -960 447498 480 0 FreeSans 448 90 0 0 la_oenb[90]
port 516 nsew signal input
flabel metal2 s 450882 -960 450994 480 0 FreeSans 448 90 0 0 la_oenb[91]
port 517 nsew signal input
flabel metal2 s 454470 -960 454582 480 0 FreeSans 448 90 0 0 la_oenb[92]
port 518 nsew signal input
flabel metal2 s 458058 -960 458170 480 0 FreeSans 448 90 0 0 la_oenb[93]
port 519 nsew signal input
flabel metal2 s 461554 -960 461666 480 0 FreeSans 448 90 0 0 la_oenb[94]
port 520 nsew signal input
flabel metal2 s 465142 -960 465254 480 0 FreeSans 448 90 0 0 la_oenb[95]
port 521 nsew signal input
flabel metal2 s 468638 -960 468750 480 0 FreeSans 448 90 0 0 la_oenb[96]
port 522 nsew signal input
flabel metal2 s 472226 -960 472338 480 0 FreeSans 448 90 0 0 la_oenb[97]
port 523 nsew signal input
flabel metal2 s 475722 -960 475834 480 0 FreeSans 448 90 0 0 la_oenb[98]
port 524 nsew signal input
flabel metal2 s 479310 -960 479422 480 0 FreeSans 448 90 0 0 la_oenb[99]
port 525 nsew signal input
flabel metal2 s 160070 -960 160182 480 0 FreeSans 448 90 0 0 la_oenb[9]
port 526 nsew signal input
flabel metal2 s 579774 -960 579886 480 0 FreeSans 448 90 0 0 user_clock2
port 527 nsew signal input
flabel metal2 s 580970 -960 581082 480 0 FreeSans 448 90 0 0 user_irq[0]
port 528 nsew signal tristate
flabel metal2 s 582166 -960 582278 480 0 FreeSans 448 90 0 0 user_irq[1]
port 529 nsew signal tristate
flabel metal2 s 583362 -960 583474 480 0 FreeSans 448 90 0 0 user_irq[2]
port 530 nsew signal tristate
flabel metal4 s -2006 -934 -1386 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 -934 585930 -314 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 704250 585930 704870 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 585310 -934 585930 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 5266 592650 5886 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 41266 592650 41886 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 77266 592650 77886 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 113266 592650 113886 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 149266 592650 149886 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 185266 592650 185886 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 221266 592650 221886 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 257266 592650 257886 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 293266 592650 293886 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 329266 592650 329886 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 365266 592650 365886 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 401266 592650 401886 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 437266 592650 437886 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 473266 592650 473886 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 509266 592650 509886 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 545266 592650 545886 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 581266 592650 581886 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 617266 592650 617886 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 653266 592650 653886 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 689266 592650 689886 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s -3926 -2854 -3306 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 -2854 587850 -2234 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 706170 587850 706790 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 587230 -2854 587850 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s -5846 -4774 -5226 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 -4774 589770 -4154 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 708090 589770 708710 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 589150 -4774 589770 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s -7766 -6694 -7146 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 -6694 591690 -6074 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 710010 591690 710630 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 591070 -6694 591690 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s -6806 -5734 -6186 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 -5734 590730 -5114 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 709050 590730 709670 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 590110 -5734 590730 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s -8726 -7654 -8106 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 -7654 592650 -7034 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 710970 592650 711590 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 592030 -7654 592650 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s -2966 -1894 -2346 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 -1894 586890 -1274 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 705210 586890 705830 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 586270 -1894 586890 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 582294 -7654 582914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 9766 592650 10386 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 45766 592650 46386 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 81766 592650 82386 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 117766 592650 118386 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 153766 592650 154386 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 189766 592650 190386 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 225766 592650 226386 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 261766 592650 262386 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 297766 592650 298386 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 333766 592650 334386 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 369766 592650 370386 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 405766 592650 406386 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 441766 592650 442386 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 477766 592650 478386 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 513766 592650 514386 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 549766 592650 550386 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 585766 592650 586386 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 621766 592650 622386 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 657766 592650 658386 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 693766 592650 694386 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s -4886 -3814 -4266 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 -3814 588810 -3194 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 707130 588810 707750 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 588190 -3814 588810 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal2 s 542 -960 654 480 0 FreeSans 448 90 0 0 wb_clk_i
port 539 nsew signal input
flabel metal2 s 1646 -960 1758 480 0 FreeSans 448 90 0 0 wb_rst_i
port 540 nsew signal input
flabel metal2 s 2842 -960 2954 480 0 FreeSans 448 90 0 0 wbs_ack_o
port 541 nsew signal tristate
flabel metal2 s 7626 -960 7738 480 0 FreeSans 448 90 0 0 wbs_adr_i[0]
port 542 nsew signal input
flabel metal2 s 47830 -960 47942 480 0 FreeSans 448 90 0 0 wbs_adr_i[10]
port 543 nsew signal input
flabel metal2 s 51326 -960 51438 480 0 FreeSans 448 90 0 0 wbs_adr_i[11]
port 544 nsew signal input
flabel metal2 s 54914 -960 55026 480 0 FreeSans 448 90 0 0 wbs_adr_i[12]
port 545 nsew signal input
flabel metal2 s 58410 -960 58522 480 0 FreeSans 448 90 0 0 wbs_adr_i[13]
port 546 nsew signal input
flabel metal2 s 61998 -960 62110 480 0 FreeSans 448 90 0 0 wbs_adr_i[14]
port 547 nsew signal input
flabel metal2 s 65494 -960 65606 480 0 FreeSans 448 90 0 0 wbs_adr_i[15]
port 548 nsew signal input
flabel metal2 s 69082 -960 69194 480 0 FreeSans 448 90 0 0 wbs_adr_i[16]
port 549 nsew signal input
flabel metal2 s 72578 -960 72690 480 0 FreeSans 448 90 0 0 wbs_adr_i[17]
port 550 nsew signal input
flabel metal2 s 76166 -960 76278 480 0 FreeSans 448 90 0 0 wbs_adr_i[18]
port 551 nsew signal input
flabel metal2 s 79662 -960 79774 480 0 FreeSans 448 90 0 0 wbs_adr_i[19]
port 552 nsew signal input
flabel metal2 s 12318 -960 12430 480 0 FreeSans 448 90 0 0 wbs_adr_i[1]
port 553 nsew signal input
flabel metal2 s 83250 -960 83362 480 0 FreeSans 448 90 0 0 wbs_adr_i[20]
port 554 nsew signal input
flabel metal2 s 86838 -960 86950 480 0 FreeSans 448 90 0 0 wbs_adr_i[21]
port 555 nsew signal input
flabel metal2 s 90334 -960 90446 480 0 FreeSans 448 90 0 0 wbs_adr_i[22]
port 556 nsew signal input
flabel metal2 s 93922 -960 94034 480 0 FreeSans 448 90 0 0 wbs_adr_i[23]
port 557 nsew signal input
flabel metal2 s 97418 -960 97530 480 0 FreeSans 448 90 0 0 wbs_adr_i[24]
port 558 nsew signal input
flabel metal2 s 101006 -960 101118 480 0 FreeSans 448 90 0 0 wbs_adr_i[25]
port 559 nsew signal input
flabel metal2 s 104502 -960 104614 480 0 FreeSans 448 90 0 0 wbs_adr_i[26]
port 560 nsew signal input
flabel metal2 s 108090 -960 108202 480 0 FreeSans 448 90 0 0 wbs_adr_i[27]
port 561 nsew signal input
flabel metal2 s 111586 -960 111698 480 0 FreeSans 448 90 0 0 wbs_adr_i[28]
port 562 nsew signal input
flabel metal2 s 115174 -960 115286 480 0 FreeSans 448 90 0 0 wbs_adr_i[29]
port 563 nsew signal input
flabel metal2 s 17010 -960 17122 480 0 FreeSans 448 90 0 0 wbs_adr_i[2]
port 564 nsew signal input
flabel metal2 s 118762 -960 118874 480 0 FreeSans 448 90 0 0 wbs_adr_i[30]
port 565 nsew signal input
flabel metal2 s 122258 -960 122370 480 0 FreeSans 448 90 0 0 wbs_adr_i[31]
port 566 nsew signal input
flabel metal2 s 21794 -960 21906 480 0 FreeSans 448 90 0 0 wbs_adr_i[3]
port 567 nsew signal input
flabel metal2 s 26486 -960 26598 480 0 FreeSans 448 90 0 0 wbs_adr_i[4]
port 568 nsew signal input
flabel metal2 s 30074 -960 30186 480 0 FreeSans 448 90 0 0 wbs_adr_i[5]
port 569 nsew signal input
flabel metal2 s 33570 -960 33682 480 0 FreeSans 448 90 0 0 wbs_adr_i[6]
port 570 nsew signal input
flabel metal2 s 37158 -960 37270 480 0 FreeSans 448 90 0 0 wbs_adr_i[7]
port 571 nsew signal input
flabel metal2 s 40654 -960 40766 480 0 FreeSans 448 90 0 0 wbs_adr_i[8]
port 572 nsew signal input
flabel metal2 s 44242 -960 44354 480 0 FreeSans 448 90 0 0 wbs_adr_i[9]
port 573 nsew signal input
flabel metal2 s 4038 -960 4150 480 0 FreeSans 448 90 0 0 wbs_cyc_i
port 574 nsew signal input
flabel metal2 s 8730 -960 8842 480 0 FreeSans 448 90 0 0 wbs_dat_i[0]
port 575 nsew signal input
flabel metal2 s 48934 -960 49046 480 0 FreeSans 448 90 0 0 wbs_dat_i[10]
port 576 nsew signal input
flabel metal2 s 52522 -960 52634 480 0 FreeSans 448 90 0 0 wbs_dat_i[11]
port 577 nsew signal input
flabel metal2 s 56018 -960 56130 480 0 FreeSans 448 90 0 0 wbs_dat_i[12]
port 578 nsew signal input
flabel metal2 s 59606 -960 59718 480 0 FreeSans 448 90 0 0 wbs_dat_i[13]
port 579 nsew signal input
flabel metal2 s 63194 -960 63306 480 0 FreeSans 448 90 0 0 wbs_dat_i[14]
port 580 nsew signal input
flabel metal2 s 66690 -960 66802 480 0 FreeSans 448 90 0 0 wbs_dat_i[15]
port 581 nsew signal input
flabel metal2 s 70278 -960 70390 480 0 FreeSans 448 90 0 0 wbs_dat_i[16]
port 582 nsew signal input
flabel metal2 s 73774 -960 73886 480 0 FreeSans 448 90 0 0 wbs_dat_i[17]
port 583 nsew signal input
flabel metal2 s 77362 -960 77474 480 0 FreeSans 448 90 0 0 wbs_dat_i[18]
port 584 nsew signal input
flabel metal2 s 80858 -960 80970 480 0 FreeSans 448 90 0 0 wbs_dat_i[19]
port 585 nsew signal input
flabel metal2 s 13514 -960 13626 480 0 FreeSans 448 90 0 0 wbs_dat_i[1]
port 586 nsew signal input
flabel metal2 s 84446 -960 84558 480 0 FreeSans 448 90 0 0 wbs_dat_i[20]
port 587 nsew signal input
flabel metal2 s 87942 -960 88054 480 0 FreeSans 448 90 0 0 wbs_dat_i[21]
port 588 nsew signal input
flabel metal2 s 91530 -960 91642 480 0 FreeSans 448 90 0 0 wbs_dat_i[22]
port 589 nsew signal input
flabel metal2 s 95118 -960 95230 480 0 FreeSans 448 90 0 0 wbs_dat_i[23]
port 590 nsew signal input
flabel metal2 s 98614 -960 98726 480 0 FreeSans 448 90 0 0 wbs_dat_i[24]
port 591 nsew signal input
flabel metal2 s 102202 -960 102314 480 0 FreeSans 448 90 0 0 wbs_dat_i[25]
port 592 nsew signal input
flabel metal2 s 105698 -960 105810 480 0 FreeSans 448 90 0 0 wbs_dat_i[26]
port 593 nsew signal input
flabel metal2 s 109286 -960 109398 480 0 FreeSans 448 90 0 0 wbs_dat_i[27]
port 594 nsew signal input
flabel metal2 s 112782 -960 112894 480 0 FreeSans 448 90 0 0 wbs_dat_i[28]
port 595 nsew signal input
flabel metal2 s 116370 -960 116482 480 0 FreeSans 448 90 0 0 wbs_dat_i[29]
port 596 nsew signal input
flabel metal2 s 18206 -960 18318 480 0 FreeSans 448 90 0 0 wbs_dat_i[2]
port 597 nsew signal input
flabel metal2 s 119866 -960 119978 480 0 FreeSans 448 90 0 0 wbs_dat_i[30]
port 598 nsew signal input
flabel metal2 s 123454 -960 123566 480 0 FreeSans 448 90 0 0 wbs_dat_i[31]
port 599 nsew signal input
flabel metal2 s 22990 -960 23102 480 0 FreeSans 448 90 0 0 wbs_dat_i[3]
port 600 nsew signal input
flabel metal2 s 27682 -960 27794 480 0 FreeSans 448 90 0 0 wbs_dat_i[4]
port 601 nsew signal input
flabel metal2 s 31270 -960 31382 480 0 FreeSans 448 90 0 0 wbs_dat_i[5]
port 602 nsew signal input
flabel metal2 s 34766 -960 34878 480 0 FreeSans 448 90 0 0 wbs_dat_i[6]
port 603 nsew signal input
flabel metal2 s 38354 -960 38466 480 0 FreeSans 448 90 0 0 wbs_dat_i[7]
port 604 nsew signal input
flabel metal2 s 41850 -960 41962 480 0 FreeSans 448 90 0 0 wbs_dat_i[8]
port 605 nsew signal input
flabel metal2 s 45438 -960 45550 480 0 FreeSans 448 90 0 0 wbs_dat_i[9]
port 606 nsew signal input
flabel metal2 s 9926 -960 10038 480 0 FreeSans 448 90 0 0 wbs_dat_o[0]
port 607 nsew signal tristate
flabel metal2 s 50130 -960 50242 480 0 FreeSans 448 90 0 0 wbs_dat_o[10]
port 608 nsew signal tristate
flabel metal2 s 53718 -960 53830 480 0 FreeSans 448 90 0 0 wbs_dat_o[11]
port 609 nsew signal tristate
flabel metal2 s 57214 -960 57326 480 0 FreeSans 448 90 0 0 wbs_dat_o[12]
port 610 nsew signal tristate
flabel metal2 s 60802 -960 60914 480 0 FreeSans 448 90 0 0 wbs_dat_o[13]
port 611 nsew signal tristate
flabel metal2 s 64298 -960 64410 480 0 FreeSans 448 90 0 0 wbs_dat_o[14]
port 612 nsew signal tristate
flabel metal2 s 67886 -960 67998 480 0 FreeSans 448 90 0 0 wbs_dat_o[15]
port 613 nsew signal tristate
flabel metal2 s 71474 -960 71586 480 0 FreeSans 448 90 0 0 wbs_dat_o[16]
port 614 nsew signal tristate
flabel metal2 s 74970 -960 75082 480 0 FreeSans 448 90 0 0 wbs_dat_o[17]
port 615 nsew signal tristate
flabel metal2 s 78558 -960 78670 480 0 FreeSans 448 90 0 0 wbs_dat_o[18]
port 616 nsew signal tristate
flabel metal2 s 82054 -960 82166 480 0 FreeSans 448 90 0 0 wbs_dat_o[19]
port 617 nsew signal tristate
flabel metal2 s 14710 -960 14822 480 0 FreeSans 448 90 0 0 wbs_dat_o[1]
port 618 nsew signal tristate
flabel metal2 s 85642 -960 85754 480 0 FreeSans 448 90 0 0 wbs_dat_o[20]
port 619 nsew signal tristate
flabel metal2 s 89138 -960 89250 480 0 FreeSans 448 90 0 0 wbs_dat_o[21]
port 620 nsew signal tristate
flabel metal2 s 92726 -960 92838 480 0 FreeSans 448 90 0 0 wbs_dat_o[22]
port 621 nsew signal tristate
flabel metal2 s 96222 -960 96334 480 0 FreeSans 448 90 0 0 wbs_dat_o[23]
port 622 nsew signal tristate
flabel metal2 s 99810 -960 99922 480 0 FreeSans 448 90 0 0 wbs_dat_o[24]
port 623 nsew signal tristate
flabel metal2 s 103306 -960 103418 480 0 FreeSans 448 90 0 0 wbs_dat_o[25]
port 624 nsew signal tristate
flabel metal2 s 106894 -960 107006 480 0 FreeSans 448 90 0 0 wbs_dat_o[26]
port 625 nsew signal tristate
flabel metal2 s 110482 -960 110594 480 0 FreeSans 448 90 0 0 wbs_dat_o[27]
port 626 nsew signal tristate
flabel metal2 s 113978 -960 114090 480 0 FreeSans 448 90 0 0 wbs_dat_o[28]
port 627 nsew signal tristate
flabel metal2 s 117566 -960 117678 480 0 FreeSans 448 90 0 0 wbs_dat_o[29]
port 628 nsew signal tristate
flabel metal2 s 19402 -960 19514 480 0 FreeSans 448 90 0 0 wbs_dat_o[2]
port 629 nsew signal tristate
flabel metal2 s 121062 -960 121174 480 0 FreeSans 448 90 0 0 wbs_dat_o[30]
port 630 nsew signal tristate
flabel metal2 s 124650 -960 124762 480 0 FreeSans 448 90 0 0 wbs_dat_o[31]
port 631 nsew signal tristate
flabel metal2 s 24186 -960 24298 480 0 FreeSans 448 90 0 0 wbs_dat_o[3]
port 632 nsew signal tristate
flabel metal2 s 28878 -960 28990 480 0 FreeSans 448 90 0 0 wbs_dat_o[4]
port 633 nsew signal tristate
flabel metal2 s 32374 -960 32486 480 0 FreeSans 448 90 0 0 wbs_dat_o[5]
port 634 nsew signal tristate
flabel metal2 s 35962 -960 36074 480 0 FreeSans 448 90 0 0 wbs_dat_o[6]
port 635 nsew signal tristate
flabel metal2 s 39550 -960 39662 480 0 FreeSans 448 90 0 0 wbs_dat_o[7]
port 636 nsew signal tristate
flabel metal2 s 43046 -960 43158 480 0 FreeSans 448 90 0 0 wbs_dat_o[8]
port 637 nsew signal tristate
flabel metal2 s 46634 -960 46746 480 0 FreeSans 448 90 0 0 wbs_dat_o[9]
port 638 nsew signal tristate
flabel metal2 s 11122 -960 11234 480 0 FreeSans 448 90 0 0 wbs_sel_i[0]
port 639 nsew signal input
flabel metal2 s 15906 -960 16018 480 0 FreeSans 448 90 0 0 wbs_sel_i[1]
port 640 nsew signal input
flabel metal2 s 20598 -960 20710 480 0 FreeSans 448 90 0 0 wbs_sel_i[2]
port 641 nsew signal input
flabel metal2 s 25290 -960 25402 480 0 FreeSans 448 90 0 0 wbs_sel_i[3]
port 642 nsew signal input
flabel metal2 s 5234 -960 5346 480 0 FreeSans 448 90 0 0 wbs_stb_i
port 643 nsew signal input
flabel metal2 s 6430 -960 6542 480 0 FreeSans 448 90 0 0 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
