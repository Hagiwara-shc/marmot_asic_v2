magic
tech sky130B
magscale 1 2
timestamp 1662338643
<< metal1 >>
rect 186498 702992 186504 703044
rect 186556 703032 186562 703044
rect 188430 703032 188436 703044
rect 186556 703004 188436 703032
rect 186556 702992 186562 703004
rect 188430 702992 188436 703004
rect 188488 702992 188494 703044
rect 235166 702992 235172 703044
rect 235224 703032 235230 703044
rect 236178 703032 236184 703044
rect 235224 703004 236184 703032
rect 235224 702992 235230 703004
rect 236178 702992 236184 703004
rect 236236 702992 236242 703044
rect 522758 702992 522764 703044
rect 522816 703032 522822 703044
rect 527082 703032 527088 703044
rect 522816 703004 527088 703032
rect 522816 702992 522822 703004
rect 527082 702992 527088 703004
rect 527140 702992 527146 703044
rect 570506 702992 570512 703044
rect 570564 703032 570570 703044
rect 575842 703032 575848 703044
rect 570564 703004 575848 703032
rect 570564 702992 570570 703004
rect 575842 702992 575848 703004
rect 575900 702992 575906 703044
rect 490926 702720 490932 702772
rect 490984 702760 490990 702772
rect 494790 702760 494796 702772
rect 490984 702732 494796 702760
rect 490984 702720 490990 702732
rect 494790 702720 494796 702732
rect 494848 702720 494854 702772
rect 538674 702720 538680 702772
rect 538732 702760 538738 702772
rect 543458 702760 543464 702772
rect 538732 702732 543464 702760
rect 538732 702720 538738 702732
rect 543458 702720 543464 702732
rect 543516 702720 543522 702772
rect 24302 702448 24308 702500
rect 24360 702488 24366 702500
rect 29270 702488 29276 702500
rect 24360 702460 29276 702488
rect 24360 702448 24366 702460
rect 29270 702448 29276 702460
rect 29328 702448 29334 702500
rect 218974 702448 218980 702500
rect 219032 702488 219038 702500
rect 220262 702488 220268 702500
rect 219032 702460 220268 702488
rect 219032 702448 219038 702460
rect 220262 702448 220268 702460
rect 220320 702448 220326 702500
rect 459094 702448 459100 702500
rect 459152 702488 459158 702500
rect 462314 702488 462320 702500
rect 459152 702460 462320 702488
rect 459152 702448 459158 702460
rect 462314 702448 462320 702460
rect 462372 702448 462378 702500
rect 506842 702448 506848 702500
rect 506900 702488 506906 702500
rect 510982 702488 510988 702500
rect 506900 702460 510988 702488
rect 506900 702448 506906 702460
rect 510982 702448 510988 702460
rect 511040 702448 511046 702500
rect 554590 702448 554596 702500
rect 554648 702488 554654 702500
rect 559650 702488 559656 702500
rect 554648 702460 559656 702488
rect 554648 702448 554654 702460
rect 559650 702448 559656 702460
rect 559708 702448 559714 702500
rect 8110 700952 8116 701004
rect 8168 700992 8174 701004
rect 13078 700992 13084 701004
rect 8168 700964 13084 700992
rect 8168 700952 8174 700964
rect 13078 700952 13084 700964
rect 13136 700952 13142 701004
rect 40494 700952 40500 701004
rect 40552 700992 40558 701004
rect 44910 700992 44916 701004
rect 40552 700964 44916 700992
rect 40552 700952 40558 700964
rect 44910 700952 44916 700964
rect 44968 700952 44974 701004
rect 56778 700952 56784 701004
rect 56836 700992 56842 701004
rect 60734 700992 60740 701004
rect 56836 700964 60740 700992
rect 56836 700952 56842 700964
rect 60734 700952 60740 700964
rect 60792 700952 60798 701004
rect 72970 700952 72976 701004
rect 73028 700992 73034 701004
rect 76742 700992 76748 701004
rect 73028 700964 76748 700992
rect 73028 700952 73034 700964
rect 76742 700952 76748 700964
rect 76800 700952 76806 701004
rect 89162 700952 89168 701004
rect 89220 700992 89226 701004
rect 92566 700992 92572 701004
rect 89220 700964 92572 700992
rect 89220 700952 89226 700964
rect 92566 700952 92572 700964
rect 92624 700952 92630 701004
rect 105446 700952 105452 701004
rect 105504 700992 105510 701004
rect 108574 700992 108580 701004
rect 105504 700964 108580 700992
rect 105504 700952 105510 700964
rect 108574 700952 108580 700964
rect 108632 700952 108638 701004
rect 121638 700952 121644 701004
rect 121696 700992 121702 701004
rect 124398 700992 124404 701004
rect 121696 700964 124404 700992
rect 121696 700952 121702 700964
rect 124398 700952 124404 700964
rect 124456 700952 124462 701004
rect 137830 700952 137836 701004
rect 137888 700992 137894 701004
rect 140406 700992 140412 701004
rect 137888 700964 140412 700992
rect 137888 700952 137894 700964
rect 140406 700952 140412 700964
rect 140464 700952 140470 701004
rect 154114 700952 154120 701004
rect 154172 700992 154178 701004
rect 156230 700992 156236 701004
rect 154172 700964 156236 700992
rect 154172 700952 154178 700964
rect 156230 700952 156236 700964
rect 156288 700952 156294 701004
rect 170306 700952 170312 701004
rect 170364 700992 170370 701004
rect 172422 700992 172428 701004
rect 170364 700964 172428 700992
rect 170364 700952 170370 700964
rect 172422 700952 172428 700964
rect 172480 700952 172486 701004
rect 202782 700952 202788 701004
rect 202840 700992 202846 701004
rect 204254 700992 204260 701004
rect 202840 700964 204260 700992
rect 202840 700952 202846 700964
rect 204254 700952 204260 700964
rect 204312 700952 204318 701004
rect 348050 700952 348056 701004
rect 348108 700992 348114 701004
rect 348786 700992 348792 701004
rect 348108 700964 348792 700992
rect 348108 700952 348114 700964
rect 348786 700952 348792 700964
rect 348844 700952 348850 701004
rect 363874 700952 363880 701004
rect 363932 700992 363938 701004
rect 364978 700992 364984 701004
rect 363932 700964 364984 700992
rect 363932 700952 363938 700964
rect 364978 700952 364984 700964
rect 365036 700952 365042 701004
rect 379330 700952 379336 701004
rect 379388 700992 379394 701004
rect 381170 700992 381176 701004
rect 379388 700964 381176 700992
rect 379388 700952 379394 700964
rect 381170 700952 381176 700964
rect 381228 700952 381234 701004
rect 395706 700952 395712 701004
rect 395764 700992 395770 701004
rect 397454 700992 397460 701004
rect 395764 700964 397460 700992
rect 395764 700952 395770 700964
rect 397454 700952 397460 700964
rect 397512 700952 397518 701004
rect 411714 700952 411720 701004
rect 411772 700992 411778 701004
rect 413646 700992 413652 701004
rect 411772 700964 413652 700992
rect 411772 700952 411778 700964
rect 413646 700952 413652 700964
rect 413704 700952 413710 701004
rect 427538 700952 427544 701004
rect 427596 700992 427602 701004
rect 429838 700992 429844 701004
rect 427596 700964 429844 700992
rect 427596 700952 427602 700964
rect 429838 700952 429844 700964
rect 429896 700952 429902 701004
rect 443546 700952 443552 701004
rect 443604 700992 443610 701004
rect 446122 700992 446128 701004
rect 443604 700964 446128 700992
rect 443604 700952 443610 700964
rect 446122 700952 446128 700964
rect 446180 700952 446186 701004
rect 475378 700952 475384 701004
rect 475436 700992 475442 701004
rect 478506 700992 478512 701004
rect 475436 700964 478512 700992
rect 475436 700952 475442 700964
rect 478506 700952 478512 700964
rect 478564 700952 478570 701004
rect 74718 3992 74724 4004
rect 60706 3964 74724 3992
rect 59722 3816 59728 3868
rect 59780 3856 59786 3868
rect 60706 3856 60734 3964
rect 74718 3952 74724 3964
rect 74776 3952 74782 4004
rect 70210 3924 70216 3936
rect 59780 3828 60734 3856
rect 61856 3896 70216 3924
rect 59780 3816 59786 3828
rect 58802 3680 58808 3732
rect 58860 3720 58866 3732
rect 61856 3720 61884 3896
rect 70210 3884 70216 3896
rect 70268 3884 70274 3936
rect 78030 3924 78036 3936
rect 76392 3896 78036 3924
rect 62022 3748 62028 3800
rect 62080 3788 62086 3800
rect 67450 3788 67456 3800
rect 62080 3760 67456 3788
rect 62080 3748 62086 3760
rect 67450 3748 67456 3760
rect 67508 3748 67514 3800
rect 76392 3788 76420 3896
rect 78030 3884 78036 3896
rect 78088 3884 78094 3936
rect 83550 3856 83556 3868
rect 67560 3760 76420 3788
rect 77496 3828 83556 3856
rect 58860 3692 61884 3720
rect 58860 3680 58866 3692
rect 63218 3612 63224 3664
rect 63276 3652 63282 3664
rect 67560 3652 67588 3760
rect 69014 3680 69020 3732
rect 69072 3720 69078 3732
rect 71406 3720 71412 3732
rect 69072 3692 71412 3720
rect 69072 3680 69078 3692
rect 71406 3680 71412 3692
rect 71464 3680 71470 3732
rect 63276 3624 67588 3652
rect 63276 3612 63282 3624
rect 69106 3612 69112 3664
rect 69164 3652 69170 3664
rect 77496 3652 77524 3828
rect 83550 3816 83556 3828
rect 83608 3816 83614 3868
rect 94590 3856 94596 3868
rect 84166 3828 94596 3856
rect 80882 3748 80888 3800
rect 80940 3788 80946 3800
rect 84166 3788 84194 3828
rect 94590 3816 94596 3828
rect 94648 3816 94654 3868
rect 122282 3816 122288 3868
rect 122340 3856 122346 3868
rect 133230 3856 133236 3868
rect 122340 3828 133236 3856
rect 122340 3816 122346 3828
rect 133230 3816 133236 3828
rect 133288 3816 133294 3868
rect 80940 3760 84194 3788
rect 80940 3748 80946 3760
rect 84470 3748 84476 3800
rect 84528 3788 84534 3800
rect 97994 3788 98000 3800
rect 84528 3760 98000 3788
rect 84528 3748 84534 3760
rect 97994 3748 98000 3760
rect 98052 3748 98058 3800
rect 114002 3748 114008 3800
rect 114060 3788 114066 3800
rect 125502 3788 125508 3800
rect 114060 3760 125508 3788
rect 114060 3748 114066 3760
rect 125502 3748 125508 3760
rect 125560 3748 125566 3800
rect 81342 3720 81348 3732
rect 69164 3624 77524 3652
rect 77588 3692 81348 3720
rect 69164 3612 69170 3624
rect 66714 3544 66720 3596
rect 66772 3584 66778 3596
rect 77588 3584 77616 3692
rect 81342 3680 81348 3692
rect 81400 3680 81406 3732
rect 85666 3680 85672 3732
rect 85724 3720 85730 3732
rect 85724 3692 87000 3720
rect 85724 3680 85730 3692
rect 86862 3652 86868 3664
rect 66772 3556 77616 3584
rect 77680 3624 86868 3652
rect 66772 3544 66778 3556
rect 56042 3476 56048 3528
rect 56100 3516 56106 3528
rect 69014 3516 69020 3528
rect 56100 3488 69020 3516
rect 56100 3476 56106 3488
rect 69014 3476 69020 3488
rect 69072 3476 69078 3528
rect 70118 3476 70124 3528
rect 70176 3516 70182 3528
rect 70176 3488 70394 3516
rect 70176 3476 70182 3488
rect 54938 3408 54944 3460
rect 54996 3448 55002 3460
rect 70210 3448 70216 3460
rect 54996 3420 70216 3448
rect 54996 3408 55002 3420
rect 70210 3408 70216 3420
rect 70268 3408 70274 3460
rect 70366 3448 70394 3488
rect 72970 3476 72976 3528
rect 73028 3516 73034 3528
rect 77680 3516 77708 3624
rect 86862 3612 86868 3624
rect 86920 3612 86926 3664
rect 86972 3652 87000 3692
rect 87782 3680 87788 3732
rect 87840 3720 87846 3732
rect 101214 3720 101220 3732
rect 87840 3692 101220 3720
rect 87840 3680 87846 3692
rect 101214 3680 101220 3692
rect 101272 3680 101278 3732
rect 116394 3680 116400 3732
rect 116452 3720 116458 3732
rect 127710 3720 127716 3732
rect 116452 3692 127716 3720
rect 116452 3680 116458 3692
rect 127710 3680 127716 3692
rect 127768 3680 127774 3732
rect 99006 3652 99012 3664
rect 86972 3624 99012 3652
rect 99006 3612 99012 3624
rect 99064 3612 99070 3664
rect 109402 3612 109408 3664
rect 109460 3652 109466 3664
rect 121178 3652 121184 3664
rect 109460 3624 121184 3652
rect 109460 3612 109466 3624
rect 121178 3612 121184 3624
rect 121236 3612 121242 3664
rect 125042 3612 125048 3664
rect 125100 3652 125106 3664
rect 135438 3652 135444 3664
rect 125100 3624 135444 3652
rect 125100 3612 125106 3624
rect 135438 3612 135444 3624
rect 135496 3612 135502 3664
rect 143626 3612 143632 3664
rect 143684 3652 143690 3664
rect 153102 3652 153108 3664
rect 143684 3624 153108 3652
rect 143684 3612 143690 3624
rect 153102 3612 153108 3624
rect 153160 3612 153166 3664
rect 82906 3584 82912 3596
rect 73028 3488 77708 3516
rect 78508 3556 82912 3584
rect 73028 3476 73034 3488
rect 78508 3448 78536 3556
rect 82906 3544 82912 3556
rect 82964 3544 82970 3596
rect 83274 3544 83280 3596
rect 83332 3584 83338 3596
rect 96798 3584 96804 3596
rect 83332 3556 96804 3584
rect 83332 3544 83338 3556
rect 96798 3544 96804 3556
rect 96856 3544 96862 3596
rect 102226 3544 102232 3596
rect 102284 3584 102290 3596
rect 114462 3584 114468 3596
rect 102284 3556 114468 3584
rect 102284 3544 102290 3556
rect 114462 3544 114468 3556
rect 114520 3544 114526 3596
rect 121086 3544 121092 3596
rect 121144 3584 121150 3596
rect 132126 3584 132132 3596
rect 121144 3556 132132 3584
rect 121144 3544 121150 3556
rect 132126 3544 132132 3556
rect 132184 3544 132190 3596
rect 136450 3544 136456 3596
rect 136508 3584 136514 3596
rect 146478 3584 146484 3596
rect 136508 3556 146484 3584
rect 136508 3544 136514 3556
rect 146478 3544 146484 3556
rect 146536 3544 146542 3596
rect 149514 3544 149520 3596
rect 149572 3584 149578 3596
rect 158622 3584 158628 3596
rect 149572 3556 158628 3584
rect 149572 3544 149578 3556
rect 158622 3544 158628 3556
rect 158680 3544 158686 3596
rect 78582 3476 78588 3528
rect 78640 3516 78646 3528
rect 92382 3516 92388 3528
rect 78640 3488 92388 3516
rect 78640 3476 78646 3488
rect 92382 3476 92388 3488
rect 92440 3476 92446 3528
rect 103606 3516 103612 3528
rect 92492 3488 103612 3516
rect 85758 3448 85764 3460
rect 70366 3420 78536 3448
rect 79428 3420 85764 3448
rect 51350 3340 51356 3392
rect 51408 3380 51414 3392
rect 66990 3380 66996 3392
rect 51408 3352 66996 3380
rect 51408 3340 51414 3352
rect 66990 3340 66996 3352
rect 67048 3340 67054 3392
rect 67450 3340 67456 3392
rect 67508 3380 67514 3392
rect 76926 3380 76932 3392
rect 67508 3352 76932 3380
rect 67508 3340 67514 3352
rect 76926 3340 76932 3352
rect 76984 3340 76990 3392
rect 65518 3272 65524 3324
rect 65576 3312 65582 3324
rect 65576 3284 70394 3312
rect 65576 3272 65582 3284
rect 50154 3204 50160 3256
rect 50212 3244 50218 3256
rect 65886 3244 65892 3256
rect 50212 3216 65892 3244
rect 50212 3204 50218 3216
rect 65886 3204 65892 3216
rect 65944 3204 65950 3256
rect 70366 3244 70394 3284
rect 71498 3272 71504 3324
rect 71556 3312 71562 3324
rect 79428 3312 79456 3420
rect 85758 3408 85764 3420
rect 85816 3408 85822 3460
rect 90358 3408 90364 3460
rect 90416 3448 90422 3460
rect 92492 3448 92520 3488
rect 103606 3476 103612 3488
rect 103664 3476 103670 3528
rect 110506 3476 110512 3528
rect 110564 3516 110570 3528
rect 122374 3516 122380 3528
rect 110564 3488 122380 3516
rect 110564 3476 110570 3488
rect 122374 3476 122380 3488
rect 122432 3476 122438 3528
rect 127066 3476 127072 3528
rect 127124 3516 127130 3528
rect 137646 3516 137652 3528
rect 127124 3488 137652 3516
rect 127124 3476 127130 3488
rect 137646 3476 137652 3488
rect 137704 3476 137710 3528
rect 139210 3476 139216 3528
rect 139268 3516 139274 3528
rect 148686 3516 148692 3528
rect 139268 3488 148692 3516
rect 139268 3476 139274 3488
rect 148686 3476 148692 3488
rect 148744 3476 148750 3528
rect 153010 3476 153016 3528
rect 153068 3516 153074 3528
rect 160186 3516 160192 3528
rect 153068 3488 160192 3516
rect 153068 3476 153074 3488
rect 160186 3476 160192 3488
rect 160244 3476 160250 3528
rect 102318 3448 102324 3460
rect 90416 3420 92520 3448
rect 93826 3420 102324 3448
rect 90416 3408 90422 3420
rect 79686 3340 79692 3392
rect 79744 3380 79750 3392
rect 82998 3380 83004 3392
rect 79744 3352 83004 3380
rect 79744 3340 79750 3352
rect 82998 3340 83004 3352
rect 83056 3340 83062 3392
rect 89530 3340 89536 3392
rect 89588 3380 89594 3392
rect 93826 3380 93854 3420
rect 102318 3408 102324 3420
rect 102376 3408 102382 3460
rect 105722 3408 105728 3460
rect 105780 3448 105786 3460
rect 117774 3448 117780 3460
rect 105780 3420 117780 3448
rect 105780 3408 105786 3420
rect 117774 3408 117780 3420
rect 117832 3408 117838 3460
rect 131758 3408 131764 3460
rect 131816 3448 131822 3460
rect 142246 3448 142252 3460
rect 131816 3420 142252 3448
rect 131816 3408 131822 3420
rect 142246 3408 142252 3420
rect 142304 3408 142310 3460
rect 142522 3408 142528 3460
rect 142580 3448 142586 3460
rect 151722 3448 151728 3460
rect 142580 3420 151728 3448
rect 142580 3408 142586 3420
rect 151722 3408 151728 3420
rect 151780 3408 151786 3460
rect 155770 3408 155776 3460
rect 155828 3448 155834 3460
rect 155828 3420 157380 3448
rect 155828 3408 155834 3420
rect 89588 3352 93854 3380
rect 89588 3340 89594 3352
rect 96246 3340 96252 3392
rect 96304 3380 96310 3392
rect 109034 3380 109040 3392
rect 96304 3352 109040 3380
rect 96304 3340 96310 3352
rect 109034 3340 109040 3352
rect 109092 3340 109098 3392
rect 112806 3340 112812 3392
rect 112864 3380 112870 3392
rect 124122 3380 124128 3392
rect 112864 3352 124128 3380
rect 112864 3340 112870 3352
rect 124122 3340 124128 3352
rect 124180 3340 124186 3392
rect 125962 3340 125968 3392
rect 126020 3380 126026 3392
rect 136634 3380 136640 3392
rect 126020 3352 136640 3380
rect 126020 3340 126026 3352
rect 136634 3340 136640 3352
rect 136692 3340 136698 3392
rect 149790 3380 149796 3392
rect 140056 3352 149796 3380
rect 71556 3284 79456 3312
rect 71556 3272 71562 3284
rect 82906 3272 82912 3324
rect 82964 3312 82970 3324
rect 84654 3312 84660 3324
rect 82964 3284 84660 3312
rect 82964 3272 82970 3284
rect 84654 3272 84660 3284
rect 84712 3272 84718 3324
rect 86862 3272 86868 3324
rect 86920 3312 86926 3324
rect 100110 3312 100116 3324
rect 86920 3284 100116 3312
rect 86920 3272 86926 3284
rect 100110 3272 100116 3284
rect 100168 3272 100174 3324
rect 103330 3272 103336 3324
rect 103388 3312 103394 3324
rect 115566 3312 115572 3324
rect 103388 3284 115572 3312
rect 103388 3272 103394 3284
rect 115566 3272 115572 3284
rect 115624 3272 115630 3324
rect 117590 3272 117596 3324
rect 117648 3312 117654 3324
rect 128814 3312 128820 3324
rect 117648 3284 128820 3312
rect 117648 3272 117654 3284
rect 128814 3272 128820 3284
rect 128872 3272 128878 3324
rect 129366 3272 129372 3324
rect 129424 3312 129430 3324
rect 139854 3312 139860 3324
rect 129424 3284 139860 3312
rect 129424 3272 129430 3284
rect 139854 3272 139860 3284
rect 139912 3272 139918 3324
rect 140056 3256 140084 3352
rect 149790 3340 149796 3352
rect 149848 3340 149854 3392
rect 148318 3272 148324 3324
rect 148376 3312 148382 3324
rect 157242 3312 157248 3324
rect 148376 3284 157248 3312
rect 148376 3272 148382 3284
rect 157242 3272 157248 3284
rect 157300 3272 157306 3324
rect 79962 3244 79968 3256
rect 70366 3216 79968 3244
rect 79962 3204 79968 3216
rect 80020 3204 80026 3256
rect 93946 3204 93952 3256
rect 94004 3244 94010 3256
rect 106734 3244 106740 3256
rect 94004 3216 106740 3244
rect 94004 3204 94010 3216
rect 106734 3204 106740 3216
rect 106792 3204 106798 3256
rect 107194 3204 107200 3256
rect 107252 3244 107258 3256
rect 118602 3244 118608 3256
rect 107252 3216 118608 3244
rect 107252 3204 107258 3216
rect 118602 3204 118608 3216
rect 118660 3204 118666 3256
rect 119890 3204 119896 3256
rect 119948 3244 119954 3256
rect 131022 3244 131028 3256
rect 119948 3216 131028 3244
rect 119948 3204 119954 3216
rect 131022 3204 131028 3216
rect 131080 3204 131086 3256
rect 140038 3204 140044 3256
rect 140096 3204 140102 3256
rect 154022 3204 154028 3256
rect 154080 3244 154086 3256
rect 154080 3216 156552 3244
rect 154080 3204 154086 3216
rect 40954 3136 40960 3188
rect 41012 3176 41018 3188
rect 57054 3176 57060 3188
rect 41012 3148 57060 3176
rect 41012 3136 41018 3148
rect 57054 3136 57060 3148
rect 57112 3136 57118 3188
rect 57514 3136 57520 3188
rect 57572 3176 57578 3188
rect 72510 3176 72516 3188
rect 57572 3148 72516 3176
rect 57572 3136 57578 3148
rect 72510 3136 72516 3148
rect 72568 3136 72574 3188
rect 73798 3136 73804 3188
rect 73856 3176 73862 3188
rect 87966 3176 87972 3188
rect 73856 3148 87972 3176
rect 73856 3136 73862 3148
rect 87966 3136 87972 3148
rect 88024 3136 88030 3188
rect 101030 3136 101036 3188
rect 101088 3176 101094 3188
rect 113082 3176 113088 3188
rect 101088 3148 113088 3176
rect 101088 3136 101094 3148
rect 113082 3136 113088 3148
rect 113140 3136 113146 3188
rect 134334 3176 134340 3188
rect 123496 3148 134340 3176
rect 52546 3068 52552 3120
rect 52604 3108 52610 3120
rect 68094 3108 68100 3120
rect 52604 3080 68100 3108
rect 52604 3068 52610 3080
rect 68094 3068 68100 3080
rect 68152 3068 68158 3120
rect 76282 3068 76288 3120
rect 76340 3108 76346 3120
rect 76340 3080 79272 3108
rect 76340 3068 76346 3080
rect 44266 3000 44272 3052
rect 44324 3040 44330 3052
rect 60366 3040 60372 3052
rect 44324 3012 60372 3040
rect 44324 3000 44330 3012
rect 60366 3000 60372 3012
rect 60424 3000 60430 3052
rect 64322 3000 64328 3052
rect 64380 3040 64386 3052
rect 79134 3040 79140 3052
rect 64380 3012 79140 3040
rect 64380 3000 64386 3012
rect 79134 3000 79140 3012
rect 79192 3000 79198 3052
rect 79244 3040 79272 3080
rect 79594 3068 79600 3120
rect 79652 3108 79658 3120
rect 89070 3108 89076 3120
rect 79652 3080 89076 3108
rect 79652 3068 79658 3080
rect 89070 3068 89076 3080
rect 89128 3068 89134 3120
rect 98730 3068 98736 3120
rect 98788 3108 98794 3120
rect 111150 3108 111156 3120
rect 98788 3080 111156 3108
rect 98788 3068 98794 3080
rect 111150 3068 111156 3080
rect 111208 3068 111214 3120
rect 111610 3068 111616 3120
rect 111668 3108 111674 3120
rect 123294 3108 123300 3120
rect 111668 3080 123300 3108
rect 111668 3068 111674 3080
rect 123294 3068 123300 3080
rect 123352 3068 123358 3120
rect 79244 3012 82860 3040
rect 33594 2932 33600 2984
rect 33652 2972 33658 2984
rect 50430 2972 50436 2984
rect 33652 2944 50436 2972
rect 33652 2932 33658 2944
rect 50430 2932 50436 2944
rect 50488 2932 50494 2984
rect 64874 2972 64880 2984
rect 50632 2944 64880 2972
rect 26602 2864 26608 2916
rect 26660 2904 26666 2916
rect 43806 2904 43812 2916
rect 26660 2876 43812 2904
rect 26660 2864 26666 2876
rect 43806 2864 43812 2876
rect 43864 2864 43870 2916
rect 48958 2864 48964 2916
rect 49016 2904 49022 2916
rect 50632 2904 50660 2944
rect 64874 2932 64880 2944
rect 64932 2932 64938 2984
rect 67910 2932 67916 2984
rect 67968 2972 67974 2984
rect 82722 2972 82728 2984
rect 67968 2944 82728 2972
rect 67968 2932 67974 2944
rect 82722 2932 82728 2944
rect 82780 2932 82786 2984
rect 82832 2972 82860 3012
rect 82998 3000 83004 3052
rect 83056 3040 83062 3052
rect 93486 3040 93492 3052
rect 83056 3012 93492 3040
rect 83056 3000 83062 3012
rect 93486 3000 93492 3012
rect 93544 3000 93550 3052
rect 95142 3000 95148 3052
rect 95200 3040 95206 3052
rect 107838 3040 107844 3052
rect 95200 3012 107844 3040
rect 95200 3000 95206 3012
rect 107838 3000 107844 3012
rect 107896 3000 107902 3052
rect 108482 3000 108488 3052
rect 108540 3040 108546 3052
rect 119982 3040 119988 3052
rect 108540 3012 119988 3040
rect 108540 3000 108546 3012
rect 119982 3000 119988 3012
rect 120040 3000 120046 3052
rect 123496 2984 123524 3148
rect 134334 3136 134340 3148
rect 134392 3136 134398 3188
rect 137646 3136 137652 3188
rect 137704 3176 137710 3188
rect 147766 3176 147772 3188
rect 137704 3148 147772 3176
rect 137704 3136 137710 3148
rect 147766 3136 147772 3148
rect 147824 3136 147830 3188
rect 156414 3176 156420 3188
rect 151556 3148 156420 3176
rect 134150 3068 134156 3120
rect 134208 3108 134214 3120
rect 144270 3108 144276 3120
rect 134208 3080 144276 3108
rect 134208 3068 134214 3080
rect 144270 3068 144276 3080
rect 144328 3068 144334 3120
rect 147122 3068 147128 3120
rect 147180 3108 147186 3120
rect 151556 3108 151584 3148
rect 156414 3136 156420 3148
rect 156472 3136 156478 3188
rect 155310 3108 155316 3120
rect 147180 3080 151584 3108
rect 151648 3080 155316 3108
rect 147180 3068 147186 3080
rect 128170 3000 128176 3052
rect 128228 3040 128234 3052
rect 138750 3040 138756 3052
rect 128228 3012 138756 3040
rect 128228 3000 128234 3012
rect 138750 3000 138756 3012
rect 138808 3000 138814 3052
rect 143166 3040 143172 3052
rect 141068 3012 143172 3040
rect 90450 2972 90456 2984
rect 82832 2944 90456 2972
rect 90450 2932 90456 2944
rect 90508 2932 90514 2984
rect 91554 2932 91560 2984
rect 91612 2972 91618 2984
rect 104526 2972 104532 2984
rect 91612 2944 104532 2972
rect 91612 2932 91618 2944
rect 104526 2932 104532 2944
rect 104584 2932 104590 2984
rect 104618 2932 104624 2984
rect 104676 2972 104682 2984
rect 116946 2972 116952 2984
rect 104676 2944 116952 2972
rect 104676 2932 104682 2944
rect 116946 2932 116952 2944
rect 117004 2932 117010 2984
rect 123478 2932 123484 2984
rect 123536 2932 123542 2984
rect 130562 2932 130568 2984
rect 130620 2972 130626 2984
rect 140958 2972 140964 2984
rect 130620 2944 140964 2972
rect 130620 2932 130626 2944
rect 140958 2932 140964 2944
rect 141016 2932 141022 2984
rect 63678 2904 63684 2916
rect 49016 2876 50660 2904
rect 55186 2876 63684 2904
rect 49016 2864 49022 2876
rect 27706 2796 27712 2848
rect 27764 2836 27770 2848
rect 45186 2836 45192 2848
rect 27764 2808 45192 2836
rect 27764 2796 27770 2808
rect 45186 2796 45192 2808
rect 45244 2796 45250 2848
rect 47854 2796 47860 2848
rect 47912 2836 47918 2848
rect 55186 2836 55214 2876
rect 63678 2864 63684 2876
rect 63736 2864 63742 2916
rect 75362 2864 75368 2916
rect 75420 2904 75426 2916
rect 79594 2904 79600 2916
rect 75420 2876 79600 2904
rect 75420 2864 75426 2876
rect 79594 2864 79600 2876
rect 79652 2864 79658 2916
rect 82078 2864 82084 2916
rect 82136 2904 82142 2916
rect 95970 2904 95976 2916
rect 82136 2876 95976 2904
rect 82136 2864 82142 2876
rect 95970 2864 95976 2876
rect 96028 2864 96034 2916
rect 97442 2864 97448 2916
rect 97500 2904 97506 2916
rect 110046 2904 110052 2916
rect 97500 2876 110052 2904
rect 97500 2864 97506 2876
rect 110046 2864 110052 2876
rect 110104 2864 110110 2916
rect 115198 2864 115204 2916
rect 115256 2904 115262 2916
rect 126882 2904 126888 2916
rect 115256 2876 126888 2904
rect 115256 2864 115262 2876
rect 126882 2864 126888 2876
rect 126940 2864 126946 2916
rect 132954 2864 132960 2916
rect 133012 2904 133018 2916
rect 141068 2904 141096 3012
rect 143166 3000 143172 3012
rect 143224 3000 143230 3052
rect 145926 3000 145932 3052
rect 145984 3040 145990 3052
rect 151648 3040 151676 3080
rect 155310 3068 155316 3080
rect 155368 3068 155374 3120
rect 156524 3108 156552 3216
rect 157352 3176 157380 3420
rect 166074 3408 166080 3460
rect 166132 3448 166138 3460
rect 166132 3420 171134 3448
rect 166132 3408 166138 3420
rect 166350 3380 166356 3392
rect 158732 3352 166356 3380
rect 158162 3272 158168 3324
rect 158220 3312 158226 3324
rect 158732 3312 158760 3352
rect 166350 3340 166356 3352
rect 166408 3340 166414 3392
rect 171106 3380 171134 3420
rect 174078 3380 174084 3392
rect 171106 3352 174084 3380
rect 174078 3340 174084 3352
rect 174136 3340 174142 3392
rect 158220 3284 158760 3312
rect 158220 3272 158226 3284
rect 161290 3272 161296 3324
rect 161348 3312 161354 3324
rect 169662 3312 169668 3324
rect 161348 3284 169668 3312
rect 161348 3272 161354 3284
rect 169662 3272 169668 3284
rect 169720 3272 169726 3324
rect 181806 3312 181812 3324
rect 174280 3284 181812 3312
rect 174280 3256 174308 3284
rect 181806 3272 181812 3284
rect 181864 3272 181870 3324
rect 564342 3272 564348 3324
rect 564400 3312 564406 3324
rect 583386 3312 583392 3324
rect 564400 3284 583392 3312
rect 564400 3272 564406 3284
rect 583386 3272 583392 3284
rect 583444 3272 583450 3324
rect 160186 3204 160192 3256
rect 160244 3244 160250 3256
rect 161934 3244 161940 3256
rect 160244 3216 161940 3244
rect 160244 3204 160250 3216
rect 161934 3204 161940 3216
rect 161992 3204 161998 3256
rect 163682 3204 163688 3256
rect 163740 3244 163746 3256
rect 171870 3244 171876 3256
rect 163740 3216 171876 3244
rect 163740 3204 163746 3216
rect 171870 3204 171876 3216
rect 171928 3204 171934 3256
rect 174262 3204 174268 3256
rect 174320 3204 174326 3256
rect 180886 3244 180892 3256
rect 178604 3216 180892 3244
rect 164142 3176 164148 3188
rect 157352 3148 164148 3176
rect 164142 3136 164148 3148
rect 164200 3136 164206 3188
rect 170766 3136 170772 3188
rect 170824 3176 170830 3188
rect 178494 3176 178500 3188
rect 170824 3148 178500 3176
rect 170824 3136 170830 3148
rect 178494 3136 178500 3148
rect 178552 3136 178558 3188
rect 162762 3108 162768 3120
rect 156524 3080 162768 3108
rect 162762 3068 162768 3080
rect 162820 3068 162826 3120
rect 164878 3068 164884 3120
rect 164936 3108 164942 3120
rect 172974 3108 172980 3120
rect 164936 3080 172980 3108
rect 164936 3068 164942 3080
rect 172974 3068 172980 3080
rect 173032 3068 173038 3120
rect 173434 3068 173440 3120
rect 173492 3108 173498 3120
rect 178604 3108 178632 3216
rect 180886 3204 180892 3216
rect 180944 3204 180950 3256
rect 184934 3204 184940 3256
rect 184992 3244 184998 3256
rect 184992 3216 190454 3244
rect 184992 3204 184998 3216
rect 181438 3136 181444 3188
rect 181496 3176 181502 3188
rect 188430 3176 188436 3188
rect 181496 3148 188436 3176
rect 181496 3136 181502 3148
rect 188430 3136 188436 3148
rect 188488 3136 188494 3188
rect 190426 3176 190454 3216
rect 200298 3204 200304 3256
rect 200356 3244 200362 3256
rect 206094 3244 206100 3256
rect 200356 3216 206100 3244
rect 200356 3204 200362 3216
rect 206094 3204 206100 3216
rect 206152 3204 206158 3256
rect 556706 3204 556712 3256
rect 556764 3244 556770 3256
rect 575106 3244 575112 3256
rect 556764 3216 575112 3244
rect 556764 3204 556770 3216
rect 575106 3204 575112 3216
rect 575164 3204 575170 3256
rect 191742 3176 191748 3188
rect 190426 3148 191748 3176
rect 191742 3136 191748 3148
rect 191800 3136 191806 3188
rect 195606 3136 195612 3188
rect 195664 3176 195670 3188
rect 201678 3176 201684 3188
rect 195664 3148 201684 3176
rect 195664 3136 195670 3148
rect 201678 3136 201684 3148
rect 201736 3136 201742 3188
rect 220262 3136 220268 3188
rect 220320 3176 220326 3188
rect 224862 3176 224868 3188
rect 220320 3148 224868 3176
rect 220320 3136 220326 3148
rect 224862 3136 224868 3148
rect 224920 3136 224926 3188
rect 561122 3136 561128 3188
rect 561180 3176 561186 3188
rect 579798 3176 579804 3188
rect 561180 3148 579804 3176
rect 561180 3136 561186 3148
rect 579798 3136 579804 3148
rect 579856 3136 579862 3188
rect 173492 3080 178632 3108
rect 173492 3068 173498 3080
rect 179046 3068 179052 3120
rect 179104 3108 179110 3120
rect 186314 3108 186320 3120
rect 179104 3080 186320 3108
rect 179104 3068 179110 3080
rect 186314 3068 186320 3080
rect 186372 3068 186378 3120
rect 190546 3068 190552 3120
rect 190604 3108 190610 3120
rect 197262 3108 197268 3120
rect 190604 3080 197268 3108
rect 190604 3068 190610 3080
rect 197262 3068 197268 3080
rect 197320 3068 197326 3120
rect 202690 3068 202696 3120
rect 202748 3108 202754 3120
rect 208302 3108 208308 3120
rect 202748 3080 208308 3108
rect 202748 3068 202754 3080
rect 208302 3068 208308 3080
rect 208360 3068 208366 3120
rect 209866 3068 209872 3120
rect 209924 3108 209930 3120
rect 214926 3108 214932 3120
rect 209924 3080 214932 3108
rect 209924 3068 209930 3080
rect 214926 3068 214932 3080
rect 214984 3068 214990 3120
rect 215662 3068 215668 3120
rect 215720 3108 215726 3120
rect 220446 3108 220452 3120
rect 215720 3080 220452 3108
rect 215720 3068 215726 3080
rect 220446 3068 220452 3080
rect 220504 3068 220510 3120
rect 221550 3068 221556 3120
rect 221608 3108 221614 3120
rect 225966 3108 225972 3120
rect 221608 3080 225972 3108
rect 221608 3068 221614 3080
rect 225966 3068 225972 3080
rect 226024 3068 226030 3120
rect 228726 3068 228732 3120
rect 228784 3108 228790 3120
rect 232590 3108 232596 3120
rect 228784 3080 232596 3108
rect 228784 3068 228790 3080
rect 232590 3068 232596 3080
rect 232648 3068 232654 3120
rect 239306 3068 239312 3120
rect 239364 3108 239370 3120
rect 242526 3108 242532 3120
rect 239364 3080 242532 3108
rect 239364 3068 239370 3080
rect 242526 3068 242532 3080
rect 242584 3068 242590 3120
rect 543458 3068 543464 3120
rect 543516 3108 543522 3120
rect 560478 3108 560484 3120
rect 543516 3080 560484 3108
rect 543516 3068 543522 3080
rect 560478 3068 560484 3080
rect 560536 3068 560542 3120
rect 562226 3068 562232 3120
rect 562284 3108 562290 3120
rect 580994 3108 581000 3120
rect 562284 3080 581000 3108
rect 562284 3068 562290 3080
rect 580994 3068 581000 3080
rect 581052 3068 581058 3120
rect 145984 3012 151676 3040
rect 145984 3000 145990 3012
rect 151814 3000 151820 3052
rect 151872 3040 151878 3052
rect 160830 3040 160836 3052
rect 151872 3012 160836 3040
rect 151872 3000 151878 3012
rect 160830 3000 160836 3012
rect 160888 3000 160894 3052
rect 162486 3000 162492 3052
rect 162544 3040 162550 3052
rect 170858 3040 170864 3052
rect 162544 3012 170864 3040
rect 162544 3000 162550 3012
rect 170858 3000 170864 3012
rect 170916 3000 170922 3052
rect 171962 3000 171968 3052
rect 172020 3040 172026 3052
rect 179598 3040 179604 3052
rect 172020 3012 179604 3040
rect 172020 3000 172026 3012
rect 179598 3000 179604 3012
rect 179656 3000 179662 3052
rect 182542 3000 182548 3052
rect 182600 3040 182606 3052
rect 189534 3040 189540 3052
rect 182600 3012 189540 3040
rect 182600 3000 182606 3012
rect 189534 3000 189540 3012
rect 189592 3000 189598 3052
rect 189718 3000 189724 3052
rect 189776 3040 189782 3052
rect 196158 3040 196164 3052
rect 189776 3012 196164 3040
rect 189776 3000 189782 3012
rect 196158 3000 196164 3012
rect 196216 3000 196222 3052
rect 200574 3040 200580 3052
rect 196360 3012 200580 3040
rect 141234 2932 141240 2984
rect 141292 2972 141298 2984
rect 150894 2972 150900 2984
rect 141292 2944 150900 2972
rect 141292 2932 141298 2944
rect 150894 2932 150900 2944
rect 150952 2932 150958 2984
rect 156598 2932 156604 2984
rect 156656 2972 156662 2984
rect 165522 2972 165528 2984
rect 156656 2944 165528 2972
rect 156656 2932 156662 2944
rect 165522 2932 165528 2944
rect 165580 2932 165586 2984
rect 167178 2932 167184 2984
rect 167236 2972 167242 2984
rect 175458 2972 175464 2984
rect 167236 2944 175464 2972
rect 167236 2932 167242 2944
rect 175458 2932 175464 2944
rect 175516 2932 175522 2984
rect 175826 2932 175832 2984
rect 175884 2972 175890 2984
rect 175884 2944 177804 2972
rect 175884 2932 175890 2944
rect 133012 2876 141096 2904
rect 133012 2864 133018 2876
rect 144730 2864 144736 2916
rect 144788 2904 144794 2916
rect 144788 2876 147674 2904
rect 144788 2864 144794 2876
rect 47912 2808 55214 2836
rect 47912 2796 47918 2808
rect 60826 2796 60832 2848
rect 60884 2836 60890 2848
rect 75822 2836 75828 2848
rect 60884 2808 75828 2836
rect 60884 2796 60890 2808
rect 75822 2796 75828 2808
rect 75880 2796 75886 2848
rect 77386 2796 77392 2848
rect 77444 2836 77450 2848
rect 91278 2836 91284 2848
rect 77444 2808 91284 2836
rect 77444 2796 77450 2808
rect 91278 2796 91284 2808
rect 91336 2796 91342 2848
rect 92750 2796 92756 2848
rect 92808 2836 92814 2848
rect 98638 2836 98644 2848
rect 92808 2808 98644 2836
rect 92808 2796 92814 2808
rect 98638 2796 98644 2808
rect 98696 2796 98702 2848
rect 99834 2796 99840 2848
rect 99892 2836 99898 2848
rect 112530 2836 112536 2848
rect 99892 2808 112536 2836
rect 99892 2796 99898 2808
rect 112530 2796 112536 2808
rect 112588 2796 112594 2848
rect 118786 2796 118792 2848
rect 118844 2836 118850 2848
rect 130194 2836 130200 2848
rect 118844 2808 130200 2836
rect 118844 2796 118850 2808
rect 130194 2796 130200 2808
rect 130252 2796 130258 2848
rect 135254 2796 135260 2848
rect 135312 2836 135318 2848
rect 145374 2836 145380 2848
rect 135312 2808 145380 2836
rect 135312 2796 135318 2808
rect 145374 2796 145380 2808
rect 145432 2796 145438 2848
rect 147646 2836 147674 2876
rect 150618 2864 150624 2916
rect 150676 2904 150682 2916
rect 160002 2904 160008 2916
rect 150676 2876 160008 2904
rect 150676 2864 150682 2876
rect 160002 2864 160008 2876
rect 160060 2864 160066 2916
rect 160094 2864 160100 2916
rect 160152 2904 160158 2916
rect 168834 2904 168840 2916
rect 160152 2876 168840 2904
rect 160152 2864 160158 2876
rect 168834 2864 168840 2876
rect 168892 2864 168898 2916
rect 169570 2864 169576 2916
rect 169628 2904 169634 2916
rect 177666 2904 177672 2916
rect 169628 2876 177672 2904
rect 169628 2864 169634 2876
rect 177666 2864 177672 2876
rect 177724 2864 177730 2916
rect 177776 2904 177804 2944
rect 177850 2932 177856 2984
rect 177908 2972 177914 2984
rect 185394 2972 185400 2984
rect 177908 2944 185400 2972
rect 177908 2932 177914 2944
rect 185394 2932 185400 2944
rect 185452 2932 185458 2984
rect 194410 2932 194416 2984
rect 194468 2972 194474 2984
rect 196360 2972 196388 3012
rect 200574 3000 200580 3012
rect 200632 3000 200638 3052
rect 203886 3000 203892 3052
rect 203944 3040 203950 3052
rect 209406 3040 209412 3052
rect 203944 3012 209412 3040
rect 203944 3000 203950 3012
rect 209406 3000 209412 3012
rect 209464 3000 209470 3052
rect 212166 3000 212172 3052
rect 212224 3040 212230 3052
rect 217134 3040 217140 3052
rect 212224 3012 217140 3040
rect 212224 3000 212230 3012
rect 217134 3000 217140 3012
rect 217192 3000 217198 3052
rect 219250 3000 219256 3052
rect 219308 3040 219314 3052
rect 223482 3040 223488 3052
rect 219308 3012 223488 3040
rect 219308 3000 219314 3012
rect 223482 3000 223488 3012
rect 223540 3000 223546 3052
rect 228174 3040 228180 3052
rect 223960 3012 228180 3040
rect 223960 2984 223988 3012
rect 228174 3000 228180 3012
rect 228232 3000 228238 3052
rect 229830 3000 229836 3052
rect 229888 3040 229894 3052
rect 233694 3040 233700 3052
rect 229888 3012 233700 3040
rect 229888 3000 229894 3012
rect 233694 3000 233700 3012
rect 233752 3000 233758 3052
rect 234614 3000 234620 3052
rect 234672 3040 234678 3052
rect 238110 3040 238116 3052
rect 234672 3012 238116 3040
rect 234672 3000 234678 3012
rect 238110 3000 238116 3012
rect 238168 3000 238174 3052
rect 240502 3000 240508 3052
rect 240560 3040 240566 3052
rect 243630 3040 243636 3052
rect 240560 3012 243636 3040
rect 240560 3000 240566 3012
rect 243630 3000 243636 3012
rect 243688 3000 243694 3052
rect 245194 3000 245200 3052
rect 245252 3040 245258 3052
rect 248046 3040 248052 3052
rect 245252 3012 248052 3040
rect 245252 3000 245258 3012
rect 248046 3000 248052 3012
rect 248104 3000 248110 3052
rect 248782 3000 248788 3052
rect 248840 3040 248846 3052
rect 251358 3040 251364 3052
rect 248840 3012 251364 3040
rect 248840 3000 248846 3012
rect 251358 3000 251364 3012
rect 251416 3000 251422 3052
rect 333698 3000 333704 3052
rect 333756 3040 333762 3052
rect 336274 3040 336280 3052
rect 333756 3012 336280 3040
rect 333756 3000 333762 3012
rect 336274 3000 336280 3012
rect 336332 3000 336338 3052
rect 530026 3000 530032 3052
rect 530084 3040 530090 3052
rect 546678 3040 546684 3052
rect 530084 3012 546684 3040
rect 530084 3000 530090 3012
rect 546678 3000 546684 3012
rect 546736 3000 546742 3052
rect 553302 3000 553308 3052
rect 553360 3040 553366 3052
rect 571518 3040 571524 3052
rect 553360 3012 571524 3040
rect 553360 3000 553366 3012
rect 571518 3000 571524 3012
rect 571576 3000 571582 3052
rect 194468 2944 196388 2972
rect 194468 2932 194474 2944
rect 199102 2932 199108 2984
rect 199160 2972 199166 2984
rect 204990 2972 204996 2984
rect 199160 2944 204996 2972
rect 199160 2932 199166 2944
rect 204990 2932 204996 2944
rect 205048 2932 205054 2984
rect 206922 2972 206928 2984
rect 205100 2944 206928 2972
rect 182910 2904 182916 2916
rect 177776 2876 182916 2904
rect 182910 2864 182916 2876
rect 182968 2864 182974 2916
rect 183738 2864 183744 2916
rect 183796 2904 183802 2916
rect 190638 2904 190644 2916
rect 183796 2876 190644 2904
rect 183796 2864 183802 2876
rect 190638 2864 190644 2876
rect 190696 2864 190702 2916
rect 192386 2864 192392 2916
rect 192444 2904 192450 2916
rect 198366 2904 198372 2916
rect 192444 2876 198372 2904
rect 192444 2864 192450 2876
rect 198366 2864 198372 2876
rect 198424 2864 198430 2916
rect 201494 2864 201500 2916
rect 201552 2904 201558 2916
rect 205100 2904 205128 2944
rect 206922 2932 206928 2944
rect 206980 2932 206986 2984
rect 208578 2932 208584 2984
rect 208636 2972 208642 2984
rect 213822 2972 213828 2984
rect 208636 2944 213828 2972
rect 208636 2932 208642 2944
rect 213822 2932 213828 2944
rect 213880 2932 213886 2984
rect 214466 2932 214472 2984
rect 214524 2972 214530 2984
rect 219342 2972 219348 2984
rect 214524 2944 219348 2972
rect 214524 2932 214530 2944
rect 219342 2932 219348 2944
rect 219400 2932 219406 2984
rect 223942 2932 223948 2984
rect 224000 2932 224006 2984
rect 225138 2932 225144 2984
rect 225196 2972 225202 2984
rect 229554 2972 229560 2984
rect 225196 2944 229560 2972
rect 225196 2932 225202 2944
rect 229554 2932 229560 2944
rect 229612 2932 229618 2984
rect 231026 2932 231032 2984
rect 231084 2972 231090 2984
rect 235074 2972 235080 2984
rect 231084 2944 235080 2972
rect 231084 2932 231090 2944
rect 235074 2932 235080 2944
rect 235132 2932 235138 2984
rect 235810 2932 235816 2984
rect 235868 2972 235874 2984
rect 239490 2972 239496 2984
rect 235868 2944 239496 2972
rect 235868 2932 235874 2944
rect 239490 2932 239496 2944
rect 239548 2932 239554 2984
rect 242066 2932 242072 2984
rect 242124 2972 242130 2984
rect 245010 2972 245016 2984
rect 242124 2944 245016 2972
rect 242124 2932 242130 2944
rect 245010 2932 245016 2944
rect 245068 2932 245074 2984
rect 247586 2932 247592 2984
rect 247644 2972 247650 2984
rect 250530 2972 250536 2984
rect 247644 2944 250536 2972
rect 247644 2932 247650 2944
rect 250530 2932 250536 2944
rect 250588 2932 250594 2984
rect 253474 2932 253480 2984
rect 253532 2972 253538 2984
rect 256050 2972 256056 2984
rect 253532 2944 256056 2972
rect 253532 2932 253538 2944
rect 256050 2932 256056 2944
rect 256108 2932 256114 2984
rect 310238 2932 310244 2984
rect 310296 2972 310302 2984
rect 311434 2972 311440 2984
rect 310296 2944 311440 2972
rect 310296 2932 310302 2944
rect 311434 2932 311440 2944
rect 311492 2932 311498 2984
rect 325694 2932 325700 2984
rect 325752 2972 325758 2984
rect 327994 2972 328000 2984
rect 325752 2944 328000 2972
rect 325752 2932 325758 2944
rect 327994 2932 328000 2944
rect 328052 2932 328058 2984
rect 329006 2932 329012 2984
rect 329064 2972 329070 2984
rect 331582 2972 331588 2984
rect 329064 2944 331588 2972
rect 329064 2932 329070 2944
rect 331582 2932 331588 2944
rect 331640 2932 331646 2984
rect 332318 2932 332324 2984
rect 332376 2972 332382 2984
rect 335078 2972 335084 2984
rect 332376 2944 335084 2972
rect 332376 2932 332382 2944
rect 335078 2932 335084 2944
rect 335136 2932 335142 2984
rect 341150 2932 341156 2984
rect 341208 2972 341214 2984
rect 344554 2972 344560 2984
rect 341208 2944 344560 2972
rect 341208 2932 341214 2944
rect 344554 2932 344560 2944
rect 344612 2932 344618 2984
rect 513282 2932 513288 2984
rect 513340 2972 513346 2984
rect 529014 2972 529020 2984
rect 513340 2944 529020 2972
rect 513340 2932 513346 2944
rect 529014 2932 529020 2944
rect 529072 2932 529078 2984
rect 549806 2932 549812 2984
rect 549864 2972 549870 2984
rect 568022 2972 568028 2984
rect 549864 2944 568028 2972
rect 549864 2932 549870 2944
rect 568022 2932 568028 2944
rect 568080 2932 568086 2984
rect 201552 2876 205128 2904
rect 201552 2864 201558 2876
rect 206186 2864 206192 2916
rect 206244 2904 206250 2916
rect 211614 2904 211620 2916
rect 206244 2876 211620 2904
rect 206244 2864 206250 2876
rect 211614 2864 211620 2876
rect 211672 2864 211678 2916
rect 213362 2864 213368 2916
rect 213420 2904 213426 2916
rect 217962 2904 217968 2916
rect 213420 2876 217968 2904
rect 213420 2864 213426 2876
rect 217962 2864 217968 2876
rect 218020 2864 218026 2916
rect 218054 2864 218060 2916
rect 218112 2904 218118 2916
rect 222930 2904 222936 2916
rect 218112 2876 222936 2904
rect 218112 2864 218118 2876
rect 222930 2864 222936 2876
rect 222988 2864 222994 2916
rect 223114 2864 223120 2916
rect 223172 2904 223178 2916
rect 227346 2904 227352 2916
rect 223172 2876 227352 2904
rect 223172 2864 223178 2876
rect 227346 2864 227352 2876
rect 227404 2864 227410 2916
rect 227530 2864 227536 2916
rect 227588 2904 227594 2916
rect 231762 2904 231768 2916
rect 227588 2876 231768 2904
rect 227588 2864 227594 2876
rect 231762 2864 231768 2876
rect 231820 2864 231826 2916
rect 232222 2864 232228 2916
rect 232280 2904 232286 2916
rect 236178 2904 236184 2916
rect 232280 2876 236184 2904
rect 232280 2864 232286 2876
rect 236178 2864 236184 2876
rect 236236 2864 236242 2916
rect 237006 2864 237012 2916
rect 237064 2904 237070 2916
rect 240594 2904 240600 2916
rect 237064 2876 240600 2904
rect 237064 2864 237070 2876
rect 240594 2864 240600 2876
rect 240652 2864 240658 2916
rect 244090 2864 244096 2916
rect 244148 2904 244154 2916
rect 247218 2904 247224 2916
rect 244148 2876 247224 2904
rect 244148 2864 244154 2876
rect 247218 2864 247224 2876
rect 247276 2864 247282 2916
rect 249978 2864 249984 2916
rect 250036 2904 250042 2916
rect 252738 2904 252744 2916
rect 250036 2876 252744 2904
rect 250036 2864 250042 2876
rect 252738 2864 252744 2876
rect 252796 2864 252802 2916
rect 254670 2864 254676 2916
rect 254728 2904 254734 2916
rect 257154 2904 257160 2916
rect 254728 2876 257160 2904
rect 254728 2864 254734 2876
rect 257154 2864 257160 2876
rect 257212 2864 257218 2916
rect 261754 2864 261760 2916
rect 261812 2904 261818 2916
rect 263778 2904 263784 2916
rect 261812 2876 263784 2904
rect 261812 2864 261818 2876
rect 263778 2864 263784 2876
rect 263836 2864 263842 2916
rect 312446 2864 312452 2916
rect 312504 2904 312510 2916
rect 313826 2904 313832 2916
rect 312504 2876 313832 2904
rect 312504 2864 312510 2876
rect 313826 2864 313832 2876
rect 313884 2864 313890 2916
rect 314562 2864 314568 2916
rect 314620 2904 314626 2916
rect 316218 2904 316224 2916
rect 314620 2876 316224 2904
rect 314620 2864 314626 2876
rect 316218 2864 316224 2876
rect 316276 2864 316282 2916
rect 316862 2864 316868 2916
rect 316920 2904 316926 2916
rect 318518 2904 318524 2916
rect 316920 2876 318524 2904
rect 316920 2864 316926 2876
rect 318518 2864 318524 2876
rect 318576 2864 318582 2916
rect 319070 2864 319076 2916
rect 319128 2904 319134 2916
rect 320910 2904 320916 2916
rect 319128 2876 320916 2904
rect 319128 2864 319134 2876
rect 320910 2864 320916 2876
rect 320968 2864 320974 2916
rect 321278 2864 321284 2916
rect 321336 2904 321342 2916
rect 323302 2904 323308 2916
rect 321336 2876 323308 2904
rect 321336 2864 321342 2876
rect 323302 2864 323308 2876
rect 323360 2864 323366 2916
rect 323486 2864 323492 2916
rect 323544 2904 323550 2916
rect 325602 2904 325608 2916
rect 323544 2876 325608 2904
rect 323544 2864 323550 2876
rect 325602 2864 325608 2876
rect 325660 2864 325666 2916
rect 327902 2864 327908 2916
rect 327960 2904 327966 2916
rect 330386 2904 330392 2916
rect 327960 2876 330392 2904
rect 327960 2864 327966 2876
rect 330386 2864 330392 2876
rect 330444 2864 330450 2916
rect 331122 2864 331128 2916
rect 331180 2904 331186 2916
rect 333882 2904 333888 2916
rect 331180 2876 333888 2904
rect 331180 2864 331186 2876
rect 333882 2864 333888 2876
rect 333940 2864 333946 2916
rect 334526 2864 334532 2916
rect 334584 2904 334590 2916
rect 337470 2904 337476 2916
rect 334584 2876 337476 2904
rect 334584 2864 334590 2876
rect 337470 2864 337476 2876
rect 337528 2864 337534 2916
rect 340046 2864 340052 2916
rect 340104 2904 340110 2916
rect 342990 2904 342996 2916
rect 340104 2876 342996 2904
rect 340104 2864 340110 2876
rect 342990 2864 342996 2876
rect 343048 2864 343054 2916
rect 517514 2864 517520 2916
rect 517572 2904 517578 2916
rect 523034 2904 523040 2916
rect 517572 2876 523040 2904
rect 517572 2864 517578 2876
rect 523034 2864 523040 2876
rect 523092 2864 523098 2916
rect 525794 2864 525800 2916
rect 525852 2904 525858 2916
rect 531314 2904 531320 2916
rect 525852 2876 531320 2904
rect 525852 2864 525858 2876
rect 531314 2864 531320 2876
rect 531372 2864 531378 2916
rect 536558 2864 536564 2916
rect 536616 2904 536622 2916
rect 553762 2904 553768 2916
rect 536616 2876 553768 2904
rect 536616 2864 536622 2876
rect 553762 2864 553768 2876
rect 553820 2864 553826 2916
rect 559742 2864 559748 2916
rect 559800 2904 559806 2916
rect 578602 2904 578608 2916
rect 559800 2876 578608 2904
rect 559800 2864 559806 2876
rect 578602 2864 578608 2876
rect 578660 2864 578666 2916
rect 154206 2836 154212 2848
rect 147646 2808 154212 2836
rect 154206 2796 154212 2808
rect 154264 2796 154270 2848
rect 158898 2796 158904 2848
rect 158956 2836 158962 2848
rect 167730 2836 167736 2848
rect 158956 2808 167736 2836
rect 158956 2796 158962 2808
rect 167730 2796 167736 2808
rect 167788 2796 167794 2848
rect 168374 2796 168380 2848
rect 168432 2836 168438 2848
rect 176286 2836 176292 2848
rect 168432 2808 176292 2836
rect 168432 2796 168438 2808
rect 176286 2796 176292 2808
rect 176344 2796 176350 2848
rect 180242 2796 180248 2848
rect 180300 2836 180306 2848
rect 187326 2836 187332 2848
rect 180300 2808 187332 2836
rect 180300 2796 180306 2808
rect 187326 2796 187332 2808
rect 187384 2796 187390 2848
rect 199470 2836 199476 2848
rect 193232 2808 199476 2836
rect 193232 2780 193260 2808
rect 199470 2796 199476 2808
rect 199528 2796 199534 2848
rect 205082 2796 205088 2848
rect 205140 2836 205146 2848
rect 210510 2836 210516 2848
rect 205140 2808 210516 2836
rect 205140 2796 205146 2808
rect 210510 2796 210516 2808
rect 210568 2796 210574 2848
rect 210970 2796 210976 2848
rect 211028 2836 211034 2848
rect 216030 2836 216036 2848
rect 211028 2808 216036 2836
rect 211028 2796 211034 2808
rect 216030 2796 216036 2808
rect 216088 2796 216094 2848
rect 216858 2796 216864 2848
rect 216916 2836 216922 2848
rect 221826 2836 221832 2848
rect 216916 2808 221832 2836
rect 216916 2796 216922 2808
rect 221826 2796 221832 2808
rect 221884 2796 221890 2848
rect 226334 2796 226340 2848
rect 226392 2836 226398 2848
rect 230658 2836 230664 2848
rect 226392 2808 230664 2836
rect 226392 2796 226398 2808
rect 230658 2796 230664 2808
rect 230716 2796 230722 2848
rect 233418 2796 233424 2848
rect 233476 2836 233482 2848
rect 237282 2836 237288 2848
rect 233476 2808 237288 2836
rect 233476 2796 233482 2808
rect 237282 2796 237288 2808
rect 237340 2796 237346 2848
rect 238110 2796 238116 2848
rect 238168 2836 238174 2848
rect 241698 2836 241704 2848
rect 238168 2808 241704 2836
rect 238168 2796 238174 2808
rect 241698 2796 241704 2808
rect 241756 2796 241762 2848
rect 242894 2796 242900 2848
rect 242952 2836 242958 2848
rect 246114 2836 246120 2848
rect 242952 2808 246120 2836
rect 242952 2796 242958 2808
rect 246114 2796 246120 2808
rect 246172 2796 246178 2848
rect 246390 2796 246396 2848
rect 246448 2836 246454 2848
rect 249426 2836 249432 2848
rect 246448 2808 249432 2836
rect 246448 2796 246454 2808
rect 249426 2796 249432 2808
rect 249484 2796 249490 2848
rect 252370 2796 252376 2848
rect 252428 2836 252434 2848
rect 254946 2836 254952 2848
rect 252428 2808 254952 2836
rect 252428 2796 252434 2808
rect 254946 2796 254952 2808
rect 255004 2796 255010 2848
rect 255866 2796 255872 2848
rect 255924 2836 255930 2848
rect 258258 2836 258264 2848
rect 255924 2808 258264 2836
rect 255924 2796 255930 2808
rect 258258 2796 258264 2808
rect 258316 2796 258322 2848
rect 260650 2796 260656 2848
rect 260708 2836 260714 2848
rect 262674 2836 262680 2848
rect 260708 2808 262680 2836
rect 260708 2796 260714 2808
rect 262674 2796 262680 2808
rect 262732 2796 262738 2848
rect 304718 2796 304724 2848
rect 304776 2836 304782 2848
rect 305546 2836 305552 2848
rect 304776 2808 305552 2836
rect 304776 2796 304782 2808
rect 305546 2796 305552 2808
rect 305604 2796 305610 2848
rect 306926 2796 306932 2848
rect 306984 2836 306990 2848
rect 307938 2836 307944 2848
rect 306984 2808 307944 2836
rect 306984 2796 306990 2808
rect 307938 2796 307944 2808
rect 307996 2796 308002 2848
rect 309134 2796 309140 2848
rect 309192 2836 309198 2848
rect 310238 2836 310244 2848
rect 309192 2808 310244 2836
rect 309192 2796 309198 2808
rect 310238 2796 310244 2808
rect 310296 2796 310302 2848
rect 311342 2796 311348 2848
rect 311400 2836 311406 2848
rect 312630 2836 312636 2848
rect 311400 2808 312636 2836
rect 311400 2796 311406 2808
rect 312630 2796 312636 2808
rect 312688 2796 312694 2848
rect 313550 2796 313556 2848
rect 313608 2836 313614 2848
rect 315022 2836 315028 2848
rect 313608 2808 315028 2836
rect 313608 2796 313614 2808
rect 315022 2796 315028 2808
rect 315080 2796 315086 2848
rect 315758 2796 315764 2848
rect 315816 2836 315822 2848
rect 317322 2836 317328 2848
rect 315816 2808 317328 2836
rect 315816 2796 315822 2808
rect 317322 2796 317328 2808
rect 317380 2796 317386 2848
rect 317966 2796 317972 2848
rect 318024 2836 318030 2848
rect 319714 2836 319720 2848
rect 318024 2808 319720 2836
rect 318024 2796 318030 2808
rect 319714 2796 319720 2808
rect 319772 2796 319778 2848
rect 320082 2796 320088 2848
rect 320140 2836 320146 2848
rect 322106 2836 322112 2848
rect 320140 2808 322112 2836
rect 320140 2796 320146 2808
rect 322106 2796 322112 2808
rect 322164 2796 322170 2848
rect 322382 2796 322388 2848
rect 322440 2836 322446 2848
rect 324406 2836 324412 2848
rect 322440 2808 324412 2836
rect 322440 2796 322446 2808
rect 324406 2796 324412 2808
rect 324464 2796 324470 2848
rect 324590 2796 324596 2848
rect 324648 2836 324654 2848
rect 326798 2836 326804 2848
rect 324648 2808 326804 2836
rect 324648 2796 324654 2808
rect 326798 2796 326804 2808
rect 326856 2796 326862 2848
rect 326982 2796 326988 2848
rect 327040 2836 327046 2848
rect 329190 2836 329196 2848
rect 327040 2808 329196 2836
rect 327040 2796 327046 2808
rect 329190 2796 329196 2808
rect 329248 2796 329254 2848
rect 330110 2796 330116 2848
rect 330168 2836 330174 2848
rect 332686 2836 332692 2848
rect 330168 2808 332692 2836
rect 330168 2796 330174 2808
rect 332686 2796 332692 2808
rect 332744 2796 332750 2848
rect 335630 2796 335636 2848
rect 335688 2836 335694 2848
rect 338666 2836 338672 2848
rect 335688 2808 338672 2836
rect 335688 2796 335694 2808
rect 338666 2796 338672 2808
rect 338724 2796 338730 2848
rect 338942 2796 338948 2848
rect 339000 2836 339006 2848
rect 342070 2836 342076 2848
rect 339000 2808 342076 2836
rect 339000 2796 339006 2808
rect 342070 2796 342076 2808
rect 342128 2796 342134 2848
rect 346670 2796 346676 2848
rect 346728 2836 346734 2848
rect 350442 2836 350448 2848
rect 346728 2808 350448 2836
rect 346728 2796 346734 2808
rect 350442 2796 350448 2808
rect 350500 2796 350506 2848
rect 353202 2796 353208 2848
rect 353260 2836 353266 2848
rect 357526 2836 357532 2848
rect 353260 2808 357532 2836
rect 353260 2796 353266 2808
rect 357526 2796 357532 2808
rect 357584 2796 357590 2848
rect 372338 2796 372344 2848
rect 372396 2836 372402 2848
rect 377674 2836 377680 2848
rect 372396 2808 377680 2836
rect 372396 2796 372402 2808
rect 377674 2796 377680 2808
rect 377732 2796 377738 2848
rect 517606 2796 517612 2848
rect 517664 2836 517670 2848
rect 521838 2836 521844 2848
rect 517664 2808 521844 2836
rect 517664 2796 517670 2808
rect 521838 2796 521844 2808
rect 521896 2796 521902 2848
rect 562962 2796 562968 2848
rect 563020 2836 563026 2848
rect 582190 2836 582196 2848
rect 563020 2808 582196 2836
rect 563020 2796 563026 2808
rect 582190 2796 582196 2808
rect 582248 2796 582254 2848
rect 193214 2728 193220 2780
rect 193272 2728 193278 2780
rect 176654 1300 176660 1352
rect 176712 1340 176718 1352
rect 184290 1340 184296 1352
rect 176712 1312 184296 1340
rect 176712 1300 176718 1312
rect 184290 1300 184296 1312
rect 184348 1300 184354 1352
rect 187326 1300 187332 1352
rect 187384 1340 187390 1352
rect 194226 1340 194232 1352
rect 187384 1312 194232 1340
rect 187384 1300 187390 1312
rect 194226 1300 194232 1312
rect 194284 1300 194290 1352
rect 198274 1300 198280 1352
rect 198332 1340 198338 1352
rect 204162 1340 204168 1352
rect 198332 1312 204168 1340
rect 198332 1300 198338 1312
rect 204162 1300 204168 1312
rect 204220 1300 204226 1352
rect 207382 1300 207388 1352
rect 207440 1340 207446 1352
rect 212994 1340 213000 1352
rect 207440 1312 213000 1340
rect 207440 1300 207446 1312
rect 212994 1300 213000 1312
rect 213052 1300 213058 1352
rect 257062 1300 257068 1352
rect 257120 1340 257126 1352
rect 259362 1340 259368 1352
rect 257120 1312 259368 1340
rect 257120 1300 257126 1312
rect 259362 1300 259368 1312
rect 259420 1300 259426 1352
rect 259454 1300 259460 1352
rect 259512 1340 259518 1352
rect 261570 1340 261576 1352
rect 259512 1312 261576 1340
rect 259512 1300 259518 1312
rect 261570 1300 261576 1312
rect 261628 1300 261634 1352
rect 262950 1300 262956 1352
rect 263008 1340 263014 1352
rect 264882 1340 264888 1352
rect 263008 1312 264888 1340
rect 263008 1300 263014 1312
rect 264882 1300 264888 1312
rect 264940 1300 264946 1352
rect 265342 1300 265348 1352
rect 265400 1340 265406 1352
rect 267090 1340 267096 1352
rect 265400 1312 267096 1340
rect 265400 1300 265406 1312
rect 267090 1300 267096 1312
rect 267148 1300 267154 1352
rect 267734 1300 267740 1352
rect 267792 1340 267798 1352
rect 269298 1340 269304 1352
rect 267792 1312 269304 1340
rect 267792 1300 267798 1312
rect 269298 1300 269304 1312
rect 269356 1300 269362 1352
rect 271230 1300 271236 1352
rect 271288 1340 271294 1352
rect 272610 1340 272616 1352
rect 271288 1312 272616 1340
rect 271288 1300 271294 1312
rect 272610 1300 272616 1312
rect 272668 1300 272674 1352
rect 273622 1300 273628 1352
rect 273680 1340 273686 1352
rect 274818 1340 274824 1352
rect 273680 1312 274824 1340
rect 273680 1300 273686 1312
rect 274818 1300 274824 1312
rect 274876 1300 274882 1352
rect 277118 1300 277124 1352
rect 277176 1340 277182 1352
rect 278130 1340 278136 1352
rect 277176 1312 278136 1340
rect 277176 1300 277182 1312
rect 278130 1300 278136 1312
rect 278188 1300 278194 1352
rect 279510 1300 279516 1352
rect 279568 1340 279574 1352
rect 280338 1340 280344 1352
rect 279568 1312 280344 1340
rect 279568 1300 279574 1312
rect 280338 1300 280344 1312
rect 280396 1300 280402 1352
rect 336642 1300 336648 1352
rect 336700 1340 336706 1352
rect 339862 1340 339868 1352
rect 336700 1312 339868 1340
rect 336700 1300 336706 1312
rect 339862 1300 339868 1312
rect 339920 1300 339926 1352
rect 342162 1300 342168 1352
rect 342220 1340 342226 1352
rect 345750 1340 345756 1352
rect 342220 1312 345756 1340
rect 342220 1300 342226 1312
rect 345750 1300 345756 1312
rect 345808 1300 345814 1352
rect 348878 1300 348884 1352
rect 348936 1340 348942 1352
rect 352834 1340 352840 1352
rect 348936 1312 352840 1340
rect 348936 1300 348942 1312
rect 352834 1300 352840 1312
rect 352892 1300 352898 1352
rect 356606 1300 356612 1352
rect 356664 1340 356670 1352
rect 361114 1340 361120 1352
rect 356664 1312 361120 1340
rect 356664 1300 356670 1312
rect 361114 1300 361120 1312
rect 361172 1300 361178 1352
rect 364242 1300 364248 1352
rect 364300 1340 364306 1352
rect 369394 1340 369400 1352
rect 364300 1312 369400 1340
rect 364300 1300 364306 1312
rect 369394 1300 369400 1312
rect 369452 1300 369458 1352
rect 374270 1300 374276 1352
rect 374328 1340 374334 1352
rect 379606 1340 379612 1352
rect 374328 1312 379612 1340
rect 374328 1300 374334 1312
rect 379606 1300 379612 1312
rect 379664 1300 379670 1352
rect 384206 1300 384212 1352
rect 384264 1340 384270 1352
rect 390646 1340 390652 1352
rect 384264 1312 390652 1340
rect 384264 1300 384270 1312
rect 390646 1300 390652 1312
rect 390704 1300 390710 1352
rect 396350 1300 396356 1352
rect 396408 1340 396414 1352
rect 403618 1340 403624 1352
rect 396408 1312 403624 1340
rect 396408 1300 396414 1312
rect 403618 1300 403624 1312
rect 403676 1300 403682 1352
rect 406286 1300 406292 1352
rect 406344 1340 406350 1352
rect 414290 1340 414296 1352
rect 406344 1312 414296 1340
rect 406344 1300 406350 1312
rect 414290 1300 414296 1312
rect 414348 1300 414354 1352
rect 419442 1300 419448 1352
rect 419500 1340 419506 1352
rect 428274 1340 428280 1352
rect 419500 1312 428280 1340
rect 419500 1300 419506 1312
rect 428274 1300 428280 1312
rect 428332 1300 428338 1352
rect 428366 1300 428372 1352
rect 428424 1340 428430 1352
rect 428424 1312 435956 1340
rect 428424 1300 428430 1312
rect 98638 1232 98644 1284
rect 98696 1272 98702 1284
rect 105906 1272 105912 1284
rect 98696 1244 105912 1272
rect 98696 1232 98702 1244
rect 105906 1232 105912 1244
rect 105964 1232 105970 1284
rect 188890 1232 188896 1284
rect 188948 1272 188954 1284
rect 195330 1272 195336 1284
rect 188948 1244 195336 1272
rect 188948 1232 188954 1244
rect 195330 1232 195336 1244
rect 195388 1232 195394 1284
rect 197170 1232 197176 1284
rect 197228 1272 197234 1284
rect 203058 1272 203064 1284
rect 197228 1244 203064 1272
rect 197228 1232 197234 1244
rect 203058 1232 203064 1244
rect 203116 1232 203122 1284
rect 258258 1232 258264 1284
rect 258316 1272 258322 1284
rect 260466 1272 260472 1284
rect 258316 1244 260472 1272
rect 258316 1232 258322 1244
rect 260466 1232 260472 1244
rect 260524 1232 260530 1284
rect 264146 1232 264152 1284
rect 264204 1272 264210 1284
rect 265986 1272 265992 1284
rect 264204 1244 265992 1272
rect 264204 1232 264210 1244
rect 265986 1232 265992 1244
rect 266044 1232 266050 1284
rect 266538 1232 266544 1284
rect 266596 1272 266602 1284
rect 268194 1272 268200 1284
rect 266596 1244 268200 1272
rect 266596 1232 266602 1244
rect 268194 1232 268200 1244
rect 268252 1232 268258 1284
rect 270034 1232 270040 1284
rect 270092 1272 270098 1284
rect 271506 1272 271512 1284
rect 270092 1244 271512 1272
rect 270092 1232 270098 1244
rect 271506 1232 271512 1244
rect 271564 1232 271570 1284
rect 272426 1232 272432 1284
rect 272484 1272 272490 1284
rect 273714 1272 273720 1284
rect 272484 1244 273720 1272
rect 272484 1232 272490 1244
rect 273714 1232 273720 1244
rect 273772 1232 273778 1284
rect 343358 1232 343364 1284
rect 343416 1272 343422 1284
rect 346946 1272 346952 1284
rect 343416 1244 346952 1272
rect 343416 1232 343422 1244
rect 346946 1232 346952 1244
rect 347004 1232 347010 1284
rect 349982 1232 349988 1284
rect 350040 1272 350046 1284
rect 354030 1272 354036 1284
rect 350040 1244 354036 1272
rect 350040 1232 350046 1244
rect 354030 1232 354036 1244
rect 354088 1232 354094 1284
rect 357710 1232 357716 1284
rect 357768 1272 357774 1284
rect 362310 1272 362316 1284
rect 357768 1244 362316 1272
rect 357768 1232 357774 1244
rect 362310 1232 362316 1244
rect 362368 1232 362374 1284
rect 365438 1232 365444 1284
rect 365496 1272 365502 1284
rect 370222 1272 370228 1284
rect 365496 1244 370228 1272
rect 365496 1232 365502 1244
rect 370222 1232 370228 1244
rect 370280 1232 370286 1284
rect 370958 1232 370964 1284
rect 371016 1272 371022 1284
rect 376110 1272 376116 1284
rect 371016 1244 376116 1272
rect 371016 1232 371022 1244
rect 376110 1232 376116 1244
rect 376168 1232 376174 1284
rect 377582 1232 377588 1284
rect 377640 1272 377646 1284
rect 383562 1272 383568 1284
rect 377640 1244 383568 1272
rect 377640 1232 377646 1244
rect 383562 1232 383568 1244
rect 383620 1232 383626 1284
rect 388622 1232 388628 1284
rect 388680 1272 388686 1284
rect 395338 1272 395344 1284
rect 388680 1244 395344 1272
rect 388680 1232 388686 1244
rect 395338 1232 395344 1244
rect 395396 1232 395402 1284
rect 404078 1232 404084 1284
rect 404136 1272 404142 1284
rect 411898 1272 411904 1284
rect 404136 1244 411904 1272
rect 404136 1232 404142 1244
rect 411898 1232 411904 1244
rect 411956 1232 411962 1284
rect 413922 1232 413928 1284
rect 413980 1272 413986 1284
rect 422570 1272 422576 1284
rect 413980 1244 422576 1272
rect 413980 1232 413986 1244
rect 422570 1232 422576 1244
rect 422628 1232 422634 1284
rect 426158 1232 426164 1284
rect 426216 1272 426222 1284
rect 435174 1272 435180 1284
rect 426216 1244 435180 1272
rect 426216 1232 426222 1244
rect 435174 1232 435180 1244
rect 435232 1232 435238 1284
rect 435928 1272 435956 1312
rect 436002 1300 436008 1352
rect 436060 1340 436066 1352
rect 436060 1312 443776 1340
rect 436060 1300 436066 1312
rect 437566 1272 437572 1284
rect 435928 1244 437572 1272
rect 437566 1232 437572 1244
rect 437624 1232 437630 1284
rect 438302 1232 438308 1284
rect 438360 1272 438366 1284
rect 443748 1272 443776 1312
rect 443822 1300 443828 1352
rect 443880 1340 443886 1352
rect 454126 1340 454132 1352
rect 443880 1312 454132 1340
rect 443880 1300 443886 1312
rect 454126 1300 454132 1312
rect 454184 1300 454190 1352
rect 456978 1340 456984 1352
rect 454788 1312 456984 1340
rect 445846 1272 445852 1284
rect 438360 1244 443684 1272
rect 443748 1244 445852 1272
rect 438360 1232 438366 1244
rect 186130 1164 186136 1216
rect 186188 1204 186194 1216
rect 193122 1204 193128 1216
rect 186188 1176 193128 1204
rect 186188 1164 186194 1176
rect 193122 1164 193128 1176
rect 193180 1164 193186 1216
rect 268838 1164 268844 1216
rect 268896 1204 268902 1216
rect 270402 1204 270408 1216
rect 268896 1176 270408 1204
rect 268896 1164 268902 1176
rect 270402 1164 270408 1176
rect 270460 1164 270466 1216
rect 359918 1164 359924 1216
rect 359976 1204 359982 1216
rect 364610 1204 364616 1216
rect 359976 1176 364616 1204
rect 359976 1164 359982 1176
rect 364610 1164 364616 1176
rect 364668 1164 364674 1216
rect 366542 1164 366548 1216
rect 366600 1204 366606 1216
rect 371326 1204 371332 1216
rect 366600 1176 371332 1204
rect 366600 1164 366606 1176
rect 371326 1164 371332 1176
rect 371384 1164 371390 1216
rect 378686 1164 378692 1216
rect 378744 1204 378750 1216
rect 384390 1204 384396 1216
rect 378744 1176 384396 1204
rect 378744 1164 378750 1176
rect 384390 1164 384396 1176
rect 384448 1164 384454 1216
rect 387518 1164 387524 1216
rect 387576 1204 387582 1216
rect 394234 1204 394240 1216
rect 387576 1176 394240 1204
rect 387576 1164 387582 1176
rect 394234 1164 394240 1176
rect 394292 1164 394298 1216
rect 395246 1164 395252 1216
rect 395304 1204 395310 1216
rect 402514 1204 402520 1216
rect 395304 1176 402520 1204
rect 395304 1164 395310 1176
rect 402514 1164 402520 1176
rect 402572 1164 402578 1216
rect 412910 1164 412916 1216
rect 412968 1204 412974 1216
rect 421374 1204 421380 1216
rect 412968 1176 421380 1204
rect 412968 1164 412974 1176
rect 421374 1164 421380 1176
rect 421432 1164 421438 1216
rect 421742 1164 421748 1216
rect 421800 1204 421806 1216
rect 430850 1204 430856 1216
rect 421800 1176 430856 1204
rect 421800 1164 421806 1176
rect 430850 1164 430856 1176
rect 430908 1164 430914 1216
rect 439406 1164 439412 1216
rect 439464 1204 439470 1216
rect 443546 1204 443552 1216
rect 439464 1176 443552 1204
rect 439464 1164 439470 1176
rect 443546 1164 443552 1176
rect 443604 1164 443610 1216
rect 443656 1204 443684 1244
rect 445846 1232 445852 1244
rect 445904 1232 445910 1284
rect 449342 1232 449348 1284
rect 449400 1272 449406 1284
rect 454788 1272 454816 1312
rect 456978 1300 456984 1312
rect 457036 1300 457042 1352
rect 457070 1300 457076 1352
rect 457128 1340 457134 1352
rect 468294 1340 468300 1352
rect 457128 1312 468300 1340
rect 457128 1300 457134 1312
rect 468294 1300 468300 1312
rect 468352 1300 468358 1352
rect 481358 1300 481364 1352
rect 481416 1340 481422 1352
rect 494698 1340 494704 1352
rect 481416 1312 494704 1340
rect 481416 1300 481422 1312
rect 494698 1300 494704 1312
rect 494756 1300 494762 1352
rect 495710 1300 495716 1352
rect 495768 1340 495774 1352
rect 509694 1340 509700 1352
rect 495768 1312 509700 1340
rect 495768 1300 495774 1312
rect 509694 1300 509700 1312
rect 509752 1300 509758 1352
rect 510062 1300 510068 1352
rect 510120 1340 510126 1352
rect 525426 1340 525432 1352
rect 510120 1312 525432 1340
rect 510120 1300 510126 1312
rect 525426 1300 525432 1312
rect 525484 1300 525490 1352
rect 539870 1300 539876 1352
rect 539928 1340 539934 1352
rect 556982 1340 556988 1352
rect 539928 1312 556988 1340
rect 539928 1300 539934 1312
rect 556982 1300 556988 1312
rect 557040 1300 557046 1352
rect 449400 1244 454816 1272
rect 449400 1232 449406 1244
rect 454862 1232 454868 1284
rect 454920 1272 454926 1284
rect 454920 1244 460934 1272
rect 454920 1232 454926 1244
rect 448606 1204 448612 1216
rect 443656 1176 448612 1204
rect 448606 1164 448612 1176
rect 448664 1164 448670 1216
rect 450446 1164 450452 1216
rect 450504 1204 450510 1216
rect 460906 1204 460934 1244
rect 462590 1232 462596 1284
rect 462648 1272 462654 1284
rect 474182 1272 474188 1284
rect 462648 1244 474188 1272
rect 462648 1232 462654 1244
rect 474182 1232 474188 1244
rect 474240 1232 474246 1284
rect 480162 1232 480168 1284
rect 480220 1272 480226 1284
rect 493134 1272 493140 1284
rect 480220 1244 493140 1272
rect 480220 1232 480226 1244
rect 493134 1232 493140 1244
rect 493192 1232 493198 1284
rect 493502 1232 493508 1284
rect 493560 1272 493566 1284
rect 507302 1272 507308 1284
rect 493560 1244 507308 1272
rect 493560 1232 493566 1244
rect 507302 1232 507308 1244
rect 507360 1232 507366 1284
rect 507762 1232 507768 1284
rect 507820 1272 507826 1284
rect 517514 1272 517520 1284
rect 507820 1244 517520 1272
rect 507820 1232 507826 1244
rect 517514 1232 517520 1244
rect 517572 1232 517578 1284
rect 534350 1232 534356 1284
rect 534408 1272 534414 1284
rect 551094 1272 551100 1284
rect 534408 1244 551100 1272
rect 534408 1232 534414 1244
rect 551094 1232 551100 1244
rect 551152 1232 551158 1284
rect 465902 1204 465908 1216
rect 450504 1176 456104 1204
rect 460906 1176 465908 1204
rect 450504 1164 450510 1176
rect 352190 1096 352196 1148
rect 352248 1136 352254 1148
rect 356330 1136 356336 1148
rect 352248 1108 356336 1136
rect 352248 1096 352254 1108
rect 356330 1096 356336 1108
rect 356388 1096 356394 1148
rect 361022 1096 361028 1148
rect 361080 1136 361086 1148
rect 365438 1136 365444 1148
rect 361080 1108 365444 1136
rect 361080 1096 361086 1108
rect 365438 1096 365444 1108
rect 365496 1096 365502 1148
rect 367646 1096 367652 1148
rect 367704 1136 367710 1148
rect 372890 1136 372896 1148
rect 367704 1108 372896 1136
rect 367704 1096 367710 1108
rect 372890 1096 372896 1108
rect 372948 1096 372954 1148
rect 375282 1096 375288 1148
rect 375340 1136 375346 1148
rect 375340 1108 379744 1136
rect 375340 1096 375346 1108
rect 4062 1028 4068 1080
rect 4120 1068 4126 1080
rect 23106 1068 23112 1080
rect 4120 1040 23112 1068
rect 4120 1028 4126 1040
rect 23106 1028 23112 1040
rect 23164 1028 23170 1080
rect 355502 1028 355508 1080
rect 355560 1068 355566 1080
rect 359918 1068 359924 1080
rect 355560 1040 359924 1068
rect 355560 1028 355566 1040
rect 359918 1028 359924 1040
rect 359976 1028 359982 1080
rect 373166 1028 373172 1080
rect 373224 1068 373230 1080
rect 378502 1068 378508 1080
rect 373224 1040 378508 1068
rect 373224 1028 373230 1040
rect 378502 1028 378508 1040
rect 378560 1028 378566 1080
rect 379716 1068 379744 1108
rect 379790 1096 379796 1148
rect 379848 1136 379854 1148
rect 385954 1136 385960 1148
rect 379848 1108 385960 1136
rect 379848 1096 379854 1108
rect 385954 1096 385960 1108
rect 386012 1096 386018 1148
rect 386322 1096 386328 1148
rect 386380 1136 386386 1148
rect 392670 1136 392676 1148
rect 386380 1108 392676 1136
rect 386380 1096 386386 1108
rect 392670 1096 392676 1108
rect 392728 1096 392734 1148
rect 397362 1096 397368 1148
rect 397420 1136 397426 1148
rect 404814 1136 404820 1148
rect 397420 1108 404820 1136
rect 397420 1096 397426 1108
rect 404814 1096 404820 1108
rect 404872 1096 404878 1148
rect 420638 1096 420644 1148
rect 420696 1136 420702 1148
rect 429286 1136 429292 1148
rect 420696 1108 429292 1136
rect 420696 1096 420702 1108
rect 429286 1096 429292 1108
rect 429344 1096 429350 1148
rect 434990 1096 434996 1148
rect 435048 1136 435054 1148
rect 445018 1136 445024 1148
rect 435048 1108 445024 1136
rect 435048 1096 435054 1108
rect 445018 1096 445024 1108
rect 445076 1096 445082 1148
rect 445202 1096 445208 1148
rect 445260 1136 445266 1148
rect 455690 1136 455696 1148
rect 445260 1108 455696 1136
rect 445260 1096 445266 1108
rect 455690 1096 455696 1108
rect 455748 1096 455754 1148
rect 456076 1136 456104 1176
rect 465902 1164 465908 1176
rect 465960 1164 465966 1216
rect 475838 1164 475844 1216
rect 475896 1204 475902 1216
rect 488810 1204 488816 1216
rect 475896 1176 488816 1204
rect 475896 1164 475902 1176
rect 488810 1164 488816 1176
rect 488868 1164 488874 1216
rect 501230 1164 501236 1216
rect 501288 1204 501294 1216
rect 515490 1204 515496 1216
rect 501288 1176 515496 1204
rect 501288 1164 501294 1176
rect 515490 1164 515496 1176
rect 515548 1164 515554 1216
rect 516686 1164 516692 1216
rect 516744 1204 516750 1216
rect 532050 1204 532056 1216
rect 516744 1176 532056 1204
rect 516744 1164 516750 1176
rect 532050 1164 532056 1176
rect 532108 1164 532114 1216
rect 461578 1136 461584 1148
rect 456076 1108 461584 1136
rect 461578 1096 461584 1108
rect 461636 1096 461642 1148
rect 469122 1096 469128 1148
rect 469180 1136 469186 1148
rect 481358 1136 481364 1148
rect 469180 1108 481364 1136
rect 469180 1096 469186 1108
rect 481358 1096 481364 1108
rect 481416 1096 481422 1148
rect 487982 1096 487988 1148
rect 488040 1136 488046 1148
rect 501414 1136 501420 1148
rect 488040 1108 501420 1136
rect 488040 1096 488046 1108
rect 501414 1096 501420 1108
rect 501472 1096 501478 1148
rect 506750 1096 506756 1148
rect 506808 1136 506814 1148
rect 517606 1136 517612 1148
rect 506808 1108 517612 1136
rect 506808 1096 506814 1108
rect 517606 1096 517612 1108
rect 517664 1096 517670 1148
rect 522206 1096 522212 1148
rect 522264 1136 522270 1148
rect 538122 1136 538128 1148
rect 522264 1108 538128 1136
rect 522264 1096 522270 1108
rect 538122 1096 538128 1108
rect 538180 1096 538186 1148
rect 381170 1068 381176 1080
rect 379716 1040 381176 1068
rect 381170 1028 381176 1040
rect 381228 1028 381234 1080
rect 385310 1028 385316 1080
rect 385368 1068 385374 1080
rect 391842 1068 391848 1080
rect 385368 1040 391848 1068
rect 385368 1028 385374 1040
rect 391842 1028 391848 1040
rect 391900 1028 391906 1080
rect 394142 1028 394148 1080
rect 394200 1068 394206 1080
rect 401318 1068 401324 1080
rect 394200 1040 401324 1068
rect 394200 1028 394206 1040
rect 401318 1028 401324 1040
rect 401376 1028 401382 1080
rect 415118 1028 415124 1080
rect 415176 1068 415182 1080
rect 423398 1068 423404 1080
rect 415176 1040 423404 1068
rect 415176 1028 415182 1040
rect 423398 1028 423404 1040
rect 423456 1028 423462 1080
rect 424962 1028 424968 1080
rect 425020 1068 425026 1080
rect 434070 1068 434076 1080
rect 425020 1040 434076 1068
rect 425020 1028 425026 1040
rect 434070 1028 434076 1040
rect 434128 1028 434134 1080
rect 441522 1028 441528 1080
rect 441580 1068 441586 1080
rect 451734 1068 451740 1080
rect 441580 1040 451740 1068
rect 441580 1028 441586 1040
rect 451734 1028 451740 1040
rect 451792 1028 451798 1080
rect 455966 1028 455972 1080
rect 456024 1068 456030 1080
rect 467466 1068 467472 1080
rect 456024 1040 467472 1068
rect 456024 1028 456030 1040
rect 467466 1028 467472 1040
rect 467524 1028 467530 1080
rect 474642 1028 474648 1080
rect 474700 1068 474706 1080
rect 487246 1068 487252 1080
rect 474700 1040 487252 1068
rect 474700 1028 474706 1040
rect 487246 1028 487252 1040
rect 487304 1028 487310 1080
rect 518802 1028 518808 1080
rect 518860 1068 518866 1080
rect 534534 1068 534540 1080
rect 518860 1040 534540 1068
rect 518860 1028 518866 1040
rect 534534 1028 534540 1040
rect 534592 1028 534598 1080
rect 20622 960 20628 1012
rect 20680 1000 20686 1012
rect 38562 1000 38568 1012
rect 20680 972 38568 1000
rect 20680 960 20686 972
rect 38562 960 38568 972
rect 38620 960 38626 1012
rect 345566 960 345572 1012
rect 345624 1000 345630 1012
rect 349246 1000 349252 1012
rect 345624 972 349252 1000
rect 345624 960 345630 972
rect 349246 960 349252 972
rect 349304 960 349310 1012
rect 351086 960 351092 1012
rect 351144 1000 351150 1012
rect 355226 1000 355232 1012
rect 351144 972 355232 1000
rect 351144 960 351150 972
rect 355226 960 355232 972
rect 355284 960 355290 1012
rect 362126 960 362132 1012
rect 362184 1000 362190 1012
rect 367002 1000 367008 1012
rect 362184 972 367008 1000
rect 362184 960 362190 972
rect 367002 960 367008 972
rect 367060 960 367066 1012
rect 369762 960 369768 1012
rect 369820 1000 369826 1012
rect 375282 1000 375288 1012
rect 369820 972 375288 1000
rect 369820 960 369826 972
rect 375282 960 375288 972
rect 375340 960 375346 1012
rect 376478 960 376484 1012
rect 376536 1000 376542 1012
rect 382366 1000 382372 1012
rect 376536 972 382372 1000
rect 376536 960 376542 972
rect 382366 960 382372 972
rect 382424 960 382430 1012
rect 422846 960 422852 1012
rect 422904 1000 422910 1012
rect 431862 1000 431868 1012
rect 422904 972 431868 1000
rect 422904 960 422910 972
rect 431862 960 431868 972
rect 431920 960 431926 1012
rect 432782 960 432788 1012
rect 432840 1000 432846 1012
rect 442626 1000 442632 1012
rect 432840 972 442632 1000
rect 432840 960 432846 972
rect 442626 960 442632 972
rect 442684 960 442690 1012
rect 443546 960 443552 1012
rect 443604 1000 443610 1012
rect 449802 1000 449808 1012
rect 443604 972 449808 1000
rect 443604 960 443610 972
rect 449802 960 449808 972
rect 449860 960 449866 1012
rect 489086 960 489092 1012
rect 489144 1000 489150 1012
rect 502978 1000 502984 1012
rect 489144 972 502984 1000
rect 489144 960 489150 972
rect 502978 960 502984 972
rect 503036 960 503042 1012
rect 519998 960 520004 1012
rect 520056 1000 520062 1012
rect 536098 1000 536104 1012
rect 520056 972 536104 1000
rect 520056 960 520062 972
rect 536098 960 536104 972
rect 536156 960 536162 1012
rect 1670 892 1676 944
rect 1728 932 1734 944
rect 20898 932 20904 944
rect 1728 904 20904 932
rect 1728 892 1734 904
rect 20898 892 20904 904
rect 20956 892 20962 944
rect 358722 892 358728 944
rect 358780 932 358786 944
rect 363506 932 363512 944
rect 358780 904 363512 932
rect 358780 892 358786 904
rect 363506 892 363512 904
rect 363564 892 363570 944
rect 416222 892 416228 944
rect 416280 932 416286 944
rect 424962 932 424968 944
rect 416280 904 424968 932
rect 416280 892 416286 904
rect 424962 892 424968 904
rect 425020 892 425026 944
rect 433886 892 433892 944
rect 433944 932 433950 944
rect 443454 932 443460 944
rect 433944 904 443460 932
rect 433944 892 433950 904
rect 443454 892 443460 904
rect 443512 892 443518 944
rect 446030 892 446036 944
rect 446088 932 446094 944
rect 456886 932 456892 944
rect 446088 904 456892 932
rect 446088 892 446094 904
rect 456886 892 456892 904
rect 456944 892 456950 944
rect 494606 892 494612 944
rect 494664 932 494670 944
rect 508866 932 508872 944
rect 494664 904 508872 932
rect 494664 892 494670 904
rect 508866 892 508872 904
rect 508924 892 508930 944
rect 515582 892 515588 944
rect 515640 932 515646 944
rect 525794 932 525800 944
rect 515640 904 525800 932
rect 515640 892 515646 904
rect 525794 892 525800 904
rect 525852 892 525858 944
rect 532142 892 532148 944
rect 532200 932 532206 944
rect 548702 932 548708 944
rect 532200 904 548708 932
rect 532200 892 532206 904
rect 548702 892 548708 904
rect 548760 892 548766 944
rect 19426 824 19432 876
rect 19484 864 19490 876
rect 37458 864 37464 876
rect 19484 836 37464 864
rect 19484 824 19490 836
rect 37458 824 37464 836
rect 37516 824 37522 876
rect 337838 824 337844 876
rect 337896 864 337902 876
rect 340966 864 340972 876
rect 337896 836 340972 864
rect 337896 824 337902 836
rect 340966 824 340972 836
rect 341024 824 341030 876
rect 347682 824 347688 876
rect 347740 864 347746 876
rect 351638 864 351644 876
rect 347740 836 351644 864
rect 347740 824 347746 836
rect 351638 824 351644 836
rect 351696 824 351702 876
rect 368750 824 368756 876
rect 368808 864 368814 876
rect 373902 864 373908 876
rect 368808 836 373908 864
rect 368808 824 368814 836
rect 373902 824 373908 836
rect 373960 824 373966 876
rect 448238 824 448244 876
rect 448296 864 448302 876
rect 459186 864 459192 876
rect 448296 836 459192 864
rect 448296 824 448302 836
rect 459186 824 459192 836
rect 459244 824 459250 876
rect 485682 824 485688 876
rect 485740 864 485746 876
rect 498930 864 498936 876
rect 485740 836 498936 864
rect 485740 824 485746 836
rect 498930 824 498936 836
rect 498988 824 498994 876
rect 527726 824 527732 876
rect 527784 864 527790 876
rect 544378 864 544384 876
rect 527784 836 544384 864
rect 527784 824 527790 836
rect 544378 824 544384 836
rect 544436 824 544442 876
rect 547598 824 547604 876
rect 547656 864 547662 876
rect 565630 864 565636 876
rect 547656 836 565636 864
rect 547656 824 547662 836
rect 565630 824 565636 836
rect 565688 824 565694 876
rect 18230 756 18236 808
rect 18288 796 18294 808
rect 36354 796 36360 808
rect 18288 768 36360 796
rect 18288 756 18294 768
rect 36354 756 36360 768
rect 36412 756 36418 808
rect 251174 756 251180 808
rect 251232 796 251238 808
rect 253842 796 253848 808
rect 251232 768 253848 796
rect 251232 756 251238 768
rect 253842 756 253848 768
rect 253900 756 253906 808
rect 427262 756 427268 808
rect 427320 796 427326 808
rect 436738 796 436744 808
rect 427320 768 436744 796
rect 427320 756 427326 768
rect 436738 756 436744 768
rect 436796 756 436802 808
rect 442718 756 442724 808
rect 442776 796 442782 808
rect 453298 796 453304 808
rect 442776 768 453304 796
rect 442776 756 442782 768
rect 453298 756 453304 768
rect 453356 756 453362 808
rect 462406 796 462412 808
rect 460906 768 462412 796
rect 9950 688 9956 740
rect 10008 728 10014 740
rect 28626 728 28632 740
rect 10008 700 28632 728
rect 10008 688 10014 700
rect 28626 688 28632 700
rect 28684 688 28690 740
rect 401870 688 401876 740
rect 401928 728 401934 740
rect 409230 728 409236 740
rect 401928 700 409236 728
rect 401928 688 401934 700
rect 409230 688 409236 700
rect 409288 688 409294 740
rect 429470 688 429476 740
rect 429528 728 429534 740
rect 439130 728 439136 740
rect 429528 700 439136 728
rect 429528 688 429534 700
rect 439130 688 439136 700
rect 439188 688 439194 740
rect 440510 688 440516 740
rect 440568 728 440574 740
rect 450906 728 450912 740
rect 440568 700 450912 728
rect 440568 688 440574 700
rect 450906 688 450912 700
rect 450964 688 450970 740
rect 451550 688 451556 740
rect 451608 728 451614 740
rect 460906 728 460934 768
rect 462406 756 462412 768
rect 462464 756 462470 808
rect 483566 756 483572 808
rect 483624 796 483630 808
rect 497090 796 497096 808
rect 483624 768 497096 796
rect 483624 756 483630 768
rect 497090 756 497096 768
rect 497148 756 497154 808
rect 499022 756 499028 808
rect 499080 796 499086 808
rect 513558 796 513564 808
rect 499080 768 513564 796
rect 499080 756 499086 768
rect 513558 756 513564 768
rect 513616 756 513622 808
rect 528830 756 528836 808
rect 528888 796 528894 808
rect 545482 796 545488 808
rect 528888 768 545488 796
rect 528888 756 528894 768
rect 545482 756 545488 768
rect 545540 756 545546 808
rect 550910 756 550916 808
rect 550968 796 550974 808
rect 569126 796 569132 808
rect 550968 768 569132 796
rect 550968 756 550974 768
rect 569126 756 569132 768
rect 569184 756 569190 808
rect 451608 700 460934 728
rect 451608 688 451614 700
rect 468110 688 468116 740
rect 468168 728 468174 740
rect 480530 728 480536 740
rect 468168 700 480536 728
rect 468168 688 468174 700
rect 480530 688 480536 700
rect 480588 688 480594 740
rect 482462 688 482468 740
rect 482520 728 482526 740
rect 495526 728 495532 740
rect 482520 700 495532 728
rect 482520 688 482526 700
rect 495526 688 495532 700
rect 495584 688 495590 740
rect 502242 688 502248 740
rect 502300 728 502306 740
rect 517146 728 517152 740
rect 502300 700 517152 728
rect 502300 688 502306 700
rect 517146 688 517152 700
rect 517204 688 517210 740
rect 521102 688 521108 740
rect 521160 728 521166 740
rect 537202 728 537208 740
rect 521160 700 537208 728
rect 521160 688 521166 700
rect 537202 688 537208 700
rect 537260 688 537266 740
rect 537662 688 537668 740
rect 537720 728 537726 740
rect 554958 728 554964 740
rect 537720 700 554964 728
rect 537720 688 537726 700
rect 554958 688 554964 700
rect 555016 688 555022 740
rect 8754 620 8760 672
rect 8812 660 8818 672
rect 27522 660 27528 672
rect 8812 632 27528 660
rect 8812 620 8818 632
rect 27522 620 27528 632
rect 27580 620 27586 672
rect 34790 620 34796 672
rect 34848 660 34854 672
rect 51810 660 51816 672
rect 34848 632 51816 660
rect 34848 620 34854 632
rect 51810 620 51816 632
rect 51868 620 51874 672
rect 393038 620 393044 672
rect 393096 660 393102 672
rect 400122 660 400128 672
rect 393096 632 400128 660
rect 393096 620 393102 632
rect 400122 620 400128 632
rect 400180 620 400186 672
rect 400766 620 400772 672
rect 400824 660 400830 672
rect 408586 660 408592 672
rect 400824 632 408592 660
rect 400824 620 400830 632
rect 408586 620 408592 632
rect 408644 620 408650 672
rect 409598 620 409604 672
rect 409656 660 409662 672
rect 417878 660 417884 672
rect 409656 632 417884 660
rect 409656 620 409662 632
rect 417878 620 417884 632
rect 417936 620 417942 672
rect 441522 660 441528 672
rect 431926 632 441528 660
rect 14734 552 14740 604
rect 14792 552 14798 604
rect 17034 552 17040 604
rect 17092 592 17098 604
rect 35250 592 35256 604
rect 17092 564 35256 592
rect 17092 552 17098 564
rect 35250 552 35256 564
rect 35308 552 35314 604
rect 35986 552 35992 604
rect 36044 592 36050 604
rect 52914 592 52920 604
rect 36044 564 52920 592
rect 36044 552 36050 564
rect 52914 552 52920 564
rect 52972 552 52978 604
rect 389726 552 389732 604
rect 389784 592 389790 604
rect 396534 592 396540 604
rect 389784 564 396540 592
rect 389784 552 389790 564
rect 396534 552 396540 564
rect 396592 552 396598 604
rect 408402 552 408408 604
rect 408460 592 408466 604
rect 416682 592 416688 604
rect 408460 564 416688 592
rect 408460 552 408466 564
rect 416682 552 416688 564
rect 416740 552 416746 604
rect 431678 552 431684 604
rect 431736 592 431742 604
rect 431926 592 431954 632
rect 441522 620 441528 632
rect 441580 620 441586 672
rect 456978 620 456984 672
rect 457036 660 457042 672
rect 460014 660 460020 672
rect 457036 632 460020 660
rect 457036 620 457042 632
rect 460014 620 460020 632
rect 460072 620 460078 672
rect 464798 620 464804 672
rect 464856 660 464862 672
rect 476942 660 476948 672
rect 464856 632 476948 660
rect 464856 620 464862 632
rect 476942 620 476948 632
rect 477000 620 477006 672
rect 486878 620 486884 672
rect 486936 660 486942 672
rect 500586 660 500592 672
rect 486936 632 500592 660
rect 486936 620 486942 632
rect 500586 620 500592 632
rect 500644 620 500650 672
rect 503438 620 503444 672
rect 503496 660 503502 672
rect 518342 660 518348 672
rect 503496 632 518348 660
rect 503496 620 503502 632
rect 518342 620 518348 632
rect 518400 620 518406 672
rect 523310 620 523316 672
rect 523368 660 523374 672
rect 523368 632 524276 660
rect 523368 620 523374 632
rect 440326 592 440332 604
rect 431736 564 431954 592
rect 438596 564 440332 592
rect 431736 552 431742 564
rect 14752 524 14780 552
rect 33042 524 33048 536
rect 14752 496 33048 524
rect 33042 484 33048 496
rect 33100 484 33106 536
rect 39758 484 39764 536
rect 39816 524 39822 536
rect 56226 524 56232 536
rect 39816 496 56232 524
rect 39816 484 39822 496
rect 56226 484 56232 496
rect 56284 484 56290 536
rect 430482 484 430488 536
rect 430540 524 430546 536
rect 438596 524 438624 564
rect 440326 552 440332 564
rect 440384 552 440390 604
rect 447042 552 447048 604
rect 447100 592 447106 604
rect 458082 592 458088 604
rect 447100 564 458088 592
rect 447100 552 447106 564
rect 458082 552 458088 564
rect 458140 552 458146 604
rect 461486 552 461492 604
rect 461544 592 461550 604
rect 473446 592 473452 604
rect 461544 564 473452 592
rect 461544 552 461550 564
rect 473446 552 473452 564
rect 473504 552 473510 604
rect 486418 552 486424 604
rect 486476 552 486482 604
rect 498194 592 498200 604
rect 489886 564 498200 592
rect 430540 496 438624 524
rect 430540 484 430546 496
rect 459462 484 459468 536
rect 459520 524 459526 536
rect 470778 524 470784 536
rect 459520 496 470784 524
rect 459520 484 459526 496
rect 470778 484 470784 496
rect 470836 484 470842 536
rect 473630 484 473636 536
rect 473688 524 473694 536
rect 486436 524 486464 552
rect 473688 496 486464 524
rect 473688 484 473694 496
rect 16206 416 16212 468
rect 16264 456 16270 468
rect 34146 456 34152 468
rect 16264 428 34152 456
rect 16264 416 16270 428
rect 34146 416 34152 428
rect 34204 416 34210 468
rect 38562 416 38568 468
rect 38620 456 38626 468
rect 55122 456 55128 468
rect 38620 428 55128 456
rect 38620 416 38626 428
rect 55122 416 55128 428
rect 55180 416 55186 468
rect 381998 416 382004 468
rect 382056 456 382062 468
rect 387886 456 387892 468
rect 382056 428 387892 456
rect 382056 416 382062 428
rect 387886 416 387892 428
rect 387944 416 387950 468
rect 412082 416 412088 468
rect 412140 456 412146 468
rect 420362 456 420368 468
rect 412140 428 420368 456
rect 412140 416 412146 428
rect 420362 416 420368 428
rect 420420 416 420426 468
rect 437198 416 437204 468
rect 437256 456 437262 468
rect 447226 456 447232 468
rect 437256 428 447232 456
rect 437256 416 437262 428
rect 447226 416 447232 428
rect 447284 416 447290 468
rect 470318 416 470324 468
rect 470376 456 470382 468
rect 482462 456 482468 468
rect 470376 428 482468 456
rect 470376 416 470382 428
rect 482462 416 482468 428
rect 482520 416 482526 468
rect 484670 416 484676 468
rect 484728 456 484734 468
rect 489886 456 489914 564
rect 498194 552 498200 564
rect 498252 552 498258 604
rect 503806 592 503812 604
rect 498396 564 503812 592
rect 484728 428 489914 456
rect 484728 416 484734 428
rect 490190 416 490196 468
rect 490248 456 490254 468
rect 498396 456 498424 564
rect 503806 552 503812 564
rect 503864 552 503870 604
rect 508958 552 508964 604
rect 509016 592 509022 604
rect 523862 592 523868 604
rect 509016 564 523868 592
rect 509016 552 509022 564
rect 523862 552 523868 564
rect 523920 552 523926 604
rect 524248 592 524276 632
rect 524322 620 524328 672
rect 524380 660 524386 672
rect 533246 660 533252 672
rect 524380 632 533252 660
rect 524380 620 524386 632
rect 533246 620 533252 632
rect 533304 620 533310 672
rect 539594 660 539600 672
rect 533356 632 539600 660
rect 533356 592 533384 632
rect 539594 620 539600 632
rect 539652 620 539658 672
rect 542078 620 542084 672
rect 542136 660 542142 672
rect 542136 632 544976 660
rect 542136 620 542142 632
rect 524248 564 533384 592
rect 533706 552 533712 604
rect 533764 552 533770 604
rect 533798 552 533804 604
rect 533856 592 533862 604
rect 533856 564 543044 592
rect 533856 552 533862 564
rect 512086 524 512092 536
rect 490248 428 498424 456
rect 499546 496 512092 524
rect 490248 416 490254 428
rect 11514 348 11520 400
rect 11572 388 11578 400
rect 29730 388 29736 400
rect 11572 360 29736 388
rect 11572 348 11578 360
rect 29730 348 29736 360
rect 29788 348 29794 400
rect 32214 348 32220 400
rect 32272 388 32278 400
rect 49602 388 49608 400
rect 32272 360 49608 388
rect 32272 348 32278 360
rect 49602 348 49608 360
rect 49660 348 49666 400
rect 407390 348 407396 400
rect 407448 388 407454 400
rect 415302 388 415308 400
rect 407448 360 415308 388
rect 407448 348 407454 360
rect 415302 348 415308 360
rect 415360 348 415366 400
rect 460566 348 460572 400
rect 460624 388 460630 400
rect 472434 388 472440 400
rect 460624 360 472440 388
rect 460624 348 460630 360
rect 472434 348 472440 360
rect 472492 348 472498 400
rect 478322 348 478328 400
rect 478380 388 478386 400
rect 490742 388 490748 400
rect 478380 360 490748 388
rect 478380 348 478386 360
rect 490742 348 490748 360
rect 490800 348 490806 400
rect 497918 348 497924 400
rect 497976 388 497982 400
rect 499546 388 499574 496
rect 512086 484 512092 496
rect 512144 484 512150 536
rect 517790 484 517796 536
rect 517848 524 517854 536
rect 533724 524 533752 552
rect 517848 496 533752 524
rect 517848 484 517854 496
rect 500126 416 500132 468
rect 500184 456 500190 468
rect 514938 456 514944 468
rect 500184 428 514944 456
rect 500184 416 500190 428
rect 514938 416 514944 428
rect 514996 416 515002 468
rect 525702 416 525708 468
rect 525760 456 525766 468
rect 542170 456 542176 468
rect 525760 428 542176 456
rect 525760 416 525766 428
rect 542170 416 542176 428
rect 542228 416 542234 468
rect 497976 360 499574 388
rect 497976 348 497982 360
rect 504542 348 504548 400
rect 504600 388 504606 400
rect 519722 388 519728 400
rect 504600 360 519728 388
rect 504600 348 504606 360
rect 519722 348 519728 360
rect 519780 348 519786 400
rect 533246 348 533252 400
rect 533304 388 533310 400
rect 540422 388 540428 400
rect 533304 360 540428 388
rect 533304 348 533310 360
rect 540422 348 540428 360
rect 540480 348 540486 400
rect 543016 388 543044 564
rect 544948 524 544976 632
rect 548978 620 548984 672
rect 549036 660 549042 672
rect 566826 660 566832 672
rect 549036 632 566832 660
rect 549036 620 549042 632
rect 566826 620 566832 632
rect 566884 620 566890 672
rect 545390 552 545396 604
rect 545448 592 545454 604
rect 563238 592 563244 604
rect 545448 564 563244 592
rect 545448 552 545454 564
rect 563238 552 563244 564
rect 563296 552 563302 604
rect 559374 524 559380 536
rect 544948 496 559380 524
rect 559374 484 559380 496
rect 559432 484 559438 536
rect 544562 416 544568 468
rect 544620 456 544626 468
rect 562226 456 562232 468
rect 544620 428 562232 456
rect 544620 416 544626 428
rect 562226 416 562232 428
rect 562284 416 562290 468
rect 550450 388 550456 400
rect 543016 360 550456 388
rect 550450 348 550456 360
rect 550508 348 550514 400
rect 555326 348 555332 400
rect 555384 388 555390 400
rect 573542 388 573548 400
rect 555384 360 573548 388
rect 555384 348 555390 360
rect 573542 348 573548 360
rect 573600 348 573606 400
rect 3234 280 3240 332
rect 3292 320 3298 332
rect 22002 320 22008 332
rect 3292 292 22008 320
rect 3292 280 3298 292
rect 22002 280 22008 292
rect 22060 280 22066 332
rect 30282 280 30288 332
rect 30340 320 30346 332
rect 47394 320 47400 332
rect 30340 292 47400 320
rect 30340 280 30346 292
rect 47394 280 47400 292
rect 47452 280 47458 332
rect 398558 280 398564 332
rect 398616 320 398622 332
rect 406194 320 406200 332
rect 398616 292 406200 320
rect 398616 280 398622 292
rect 406194 280 406200 292
rect 406252 280 406258 332
rect 410978 280 410984 332
rect 411036 320 411042 332
rect 418614 320 418620 332
rect 411036 292 418620 320
rect 411036 280 411042 292
rect 418614 280 418620 292
rect 418672 280 418678 332
rect 453758 280 453764 332
rect 453816 320 453822 332
rect 464982 320 464988 332
rect 453816 292 464988 320
rect 453816 280 453822 292
rect 464982 280 464988 292
rect 465040 280 465046 332
rect 471422 280 471428 332
rect 471480 320 471486 332
rect 484210 320 484216 332
rect 471480 292 484216 320
rect 471480 280 471486 292
rect 484210 280 484216 292
rect 484268 280 484274 332
rect 505646 280 505652 332
rect 505704 320 505710 332
rect 520366 320 520372 332
rect 505704 292 520372 320
rect 505704 280 505710 292
rect 520366 280 520372 292
rect 520424 280 520430 332
rect 531038 280 531044 332
rect 531096 320 531102 332
rect 548058 320 548064 332
rect 531096 292 548064 320
rect 531096 280 531102 292
rect 548058 280 548064 292
rect 548116 280 548122 332
rect 551922 280 551928 332
rect 551980 320 551986 332
rect 570506 320 570512 332
rect 551980 292 570512 320
rect 551980 280 551986 292
rect 570506 280 570512 292
rect 570564 280 570570 332
rect 22830 212 22836 264
rect 22888 252 22894 264
rect 40494 252 40500 264
rect 22888 224 40500 252
rect 22888 212 22894 224
rect 40494 212 40500 224
rect 40552 212 40558 264
rect 42242 212 42248 264
rect 42300 252 42306 264
rect 58158 252 58164 264
rect 42300 224 58164 252
rect 42300 212 42306 224
rect 58158 212 58164 224
rect 58216 212 58222 264
rect 354398 212 354404 264
rect 354456 252 354462 264
rect 358906 252 358912 264
rect 354456 224 358912 252
rect 354456 212 354462 224
rect 358906 212 358912 224
rect 358964 212 358970 264
rect 380802 212 380808 264
rect 380860 252 380866 264
rect 386782 252 386788 264
rect 380860 224 386788 252
rect 380860 212 380866 224
rect 386782 212 386788 224
rect 386840 212 386846 264
rect 391658 212 391664 264
rect 391716 252 391722 264
rect 398742 252 398748 264
rect 391716 224 398748 252
rect 391716 212 391722 224
rect 398742 212 398748 224
rect 398800 212 398806 264
rect 405182 212 405188 264
rect 405240 252 405246 264
rect 412818 252 412824 264
rect 405240 224 412824 252
rect 405240 212 405246 224
rect 412818 212 412824 224
rect 412876 212 412882 264
rect 457898 212 457904 264
rect 457956 252 457962 264
rect 470042 252 470048 264
rect 457956 224 470048 252
rect 457956 212 457962 224
rect 470042 212 470048 224
rect 470100 212 470106 264
rect 472526 212 472532 264
rect 472584 252 472590 264
rect 484854 252 484860 264
rect 472584 224 484860 252
rect 472584 212 472590 224
rect 484854 212 484860 224
rect 484912 212 484918 264
rect 511442 212 511448 264
rect 511500 252 511506 264
rect 526254 252 526260 264
rect 511500 224 526260 252
rect 511500 212 511506 224
rect 526254 212 526260 224
rect 526312 212 526318 264
rect 538766 212 538772 264
rect 538824 252 538830 264
rect 556338 252 556344 264
rect 538824 224 556344 252
rect 538824 212 538830 224
rect 556338 212 556344 224
rect 556396 212 556402 264
rect 557166 212 557172 264
rect 557224 252 557230 264
rect 575934 252 575940 264
rect 557224 224 575940 252
rect 557224 212 557230 224
rect 575934 212 575940 224
rect 575992 212 575998 264
rect 8018 144 8024 196
rect 8076 184 8082 196
rect 26326 184 26332 196
rect 8076 156 26332 184
rect 8076 144 8082 156
rect 26326 144 26332 156
rect 26384 144 26390 196
rect 31110 144 31116 196
rect 31168 184 31174 196
rect 48498 184 48504 196
rect 31168 156 48504 184
rect 31168 144 31174 156
rect 48498 144 48504 156
rect 48556 144 48562 196
rect 53558 144 53564 196
rect 53616 184 53622 196
rect 69474 184 69480 196
rect 53616 156 69480 184
rect 53616 144 53622 156
rect 69474 144 69480 156
rect 69532 144 69538 196
rect 418430 144 418436 196
rect 418488 184 418494 196
rect 426894 184 426900 196
rect 418488 156 426900 184
rect 418488 144 418494 156
rect 426894 144 426900 156
rect 426952 144 426958 196
rect 465810 144 465816 196
rect 465868 184 465874 196
rect 478322 184 478328 196
rect 465868 156 478328 184
rect 465868 144 465874 156
rect 478322 144 478328 156
rect 478380 144 478386 196
rect 479150 144 479156 196
rect 479208 184 479214 196
rect 492490 184 492496 196
rect 479208 156 492496 184
rect 479208 144 479214 156
rect 492490 144 492496 156
rect 492548 144 492554 196
rect 492582 144 492588 196
rect 492640 184 492646 196
rect 506658 184 506664 196
rect 492640 156 506664 184
rect 492640 144 492646 156
rect 506658 144 506664 156
rect 506716 144 506722 196
rect 512638 144 512644 196
rect 512696 184 512702 196
rect 528002 184 528008 196
rect 512696 156 528008 184
rect 512696 144 512702 156
rect 528002 144 528008 156
rect 528060 144 528066 196
rect 535362 144 535368 196
rect 535420 184 535426 196
rect 552842 184 552848 196
rect 535420 156 552848 184
rect 535420 144 535426 156
rect 552842 144 552848 156
rect 552900 144 552906 196
rect 554222 144 554228 196
rect 554280 184 554286 196
rect 572898 184 572904 196
rect 554280 156 572904 184
rect 554280 144 554286 156
rect 572898 144 572904 156
rect 572956 144 572962 196
rect 22002 76 22008 128
rect 22060 116 22066 128
rect 39390 116 39396 128
rect 22060 88 39396 116
rect 22060 76 22066 88
rect 39390 76 39396 88
rect 39448 76 39454 128
rect 45278 76 45284 128
rect 45336 116 45342 128
rect 61746 116 61752 128
rect 45336 88 61752 116
rect 45336 76 45342 88
rect 61746 76 61752 88
rect 61804 76 61810 128
rect 399662 76 399668 128
rect 399720 116 399726 128
rect 407022 116 407028 128
rect 399720 88 407028 116
rect 399720 76 399726 88
rect 407022 76 407028 88
rect 407080 76 407086 128
rect 423950 76 423956 128
rect 424008 116 424014 128
rect 433426 116 433432 128
rect 424008 88 433432 116
rect 424008 76 424014 88
rect 433426 76 433432 88
rect 433484 76 433490 128
rect 452562 76 452568 128
rect 452620 116 452626 128
rect 464154 116 464160 128
rect 452620 88 464160 116
rect 452620 76 452626 88
rect 464154 76 464160 88
rect 464212 76 464218 128
rect 467006 76 467012 128
rect 467064 116 467070 128
rect 478966 116 478972 128
rect 467064 88 478972 116
rect 467064 76 467070 88
rect 478966 76 478972 88
rect 479024 76 479030 128
rect 491294 76 491300 128
rect 491352 116 491358 128
rect 505554 116 505560 128
rect 491352 88 505560 116
rect 491352 76 491358 88
rect 505554 76 505560 88
rect 505612 76 505618 128
rect 514478 76 514484 128
rect 514536 116 514542 128
rect 529934 116 529940 128
rect 514536 88 529940 116
rect 514536 76 514542 88
rect 529934 76 529940 88
rect 529992 76 529998 128
rect 540974 76 540980 128
rect 541032 116 541038 128
rect 558730 116 558736 128
rect 541032 88 558736 116
rect 541032 76 541038 88
rect 558730 76 558736 88
rect 558788 76 558794 128
rect 558822 76 558828 128
rect 558880 116 558886 128
rect 577130 116 577136 128
rect 558880 88 577136 116
rect 558880 76 558886 88
rect 577130 76 577136 88
rect 577188 76 577194 128
rect 382 8 388 60
rect 440 48 446 60
rect 19794 48 19800 60
rect 440 20 19800 48
rect 440 8 446 20
rect 19794 8 19800 20
rect 19852 8 19858 60
rect 24578 8 24584 60
rect 24636 48 24642 60
rect 41598 48 41604 60
rect 24636 20 41604 48
rect 24636 8 24642 20
rect 41598 8 41604 20
rect 41656 8 41662 60
rect 42886 8 42892 60
rect 42944 48 42950 60
rect 59354 48 59360 60
rect 42944 20 59360 48
rect 42944 8 42950 20
rect 59354 8 59360 20
rect 59412 8 59418 60
rect 344738 8 344744 60
rect 344796 48 344802 60
rect 348234 48 348240 60
rect 344796 20 348240 48
rect 344796 8 344802 20
rect 348234 8 348240 20
rect 348292 8 348298 60
rect 363230 8 363236 60
rect 363288 48 363294 60
rect 367830 48 367836 60
rect 363288 20 367836 48
rect 363288 8 363294 20
rect 367830 8 367836 20
rect 367888 8 367894 60
rect 383102 8 383108 60
rect 383160 48 383166 60
rect 389634 48 389640 60
rect 383160 20 389640 48
rect 383160 8 383166 20
rect 389634 8 389640 20
rect 389692 8 389698 60
rect 390830 8 390836 60
rect 390888 48 390894 60
rect 397914 48 397920 60
rect 390888 20 397920 48
rect 390888 8 390894 20
rect 397914 8 397920 20
rect 397972 8 397978 60
rect 402882 8 402888 60
rect 402940 48 402946 60
rect 410978 48 410984 60
rect 402940 20 410984 48
rect 402940 8 402946 20
rect 410978 8 410984 20
rect 411036 8 411042 60
rect 417326 8 417332 60
rect 417384 48 417390 60
rect 425790 48 425796 60
rect 417384 20 425796 48
rect 417384 8 417390 20
rect 425790 8 425796 20
rect 425848 8 425854 60
rect 463602 8 463608 60
rect 463660 48 463666 60
rect 475930 48 475936 60
rect 463660 20 475936 48
rect 463660 8 463666 20
rect 475930 8 475936 20
rect 475988 8 475994 60
rect 477218 8 477224 60
rect 477276 48 477282 60
rect 490098 48 490104 60
rect 477276 20 490104 48
rect 477276 8 477282 20
rect 490098 8 490104 20
rect 490156 8 490162 60
rect 496722 8 496728 60
rect 496780 48 496786 60
rect 511442 48 511448 60
rect 496780 20 511448 48
rect 496780 8 496786 20
rect 511442 8 511448 20
rect 511500 8 511506 60
rect 526898 8 526904 60
rect 526956 48 526962 60
rect 542814 48 542820 60
rect 526956 20 542820 48
rect 526956 8 526962 20
rect 542814 8 542820 20
rect 542872 8 542878 60
rect 546402 8 546408 60
rect 546460 48 546466 60
rect 564618 48 564624 60
rect 546460 20 564624 48
rect 546460 8 546466 20
rect 564618 8 564624 20
rect 564676 8 564682 60
<< via1 >>
rect 186504 702992 186556 703044
rect 188436 702992 188488 703044
rect 235172 702992 235224 703044
rect 236184 702992 236236 703044
rect 522764 702992 522816 703044
rect 527088 702992 527140 703044
rect 570512 702992 570564 703044
rect 575848 702992 575900 703044
rect 490932 702720 490984 702772
rect 494796 702720 494848 702772
rect 538680 702720 538732 702772
rect 543464 702720 543516 702772
rect 24308 702448 24360 702500
rect 29276 702448 29328 702500
rect 218980 702448 219032 702500
rect 220268 702448 220320 702500
rect 459100 702448 459152 702500
rect 462320 702448 462372 702500
rect 506848 702448 506900 702500
rect 510988 702448 511040 702500
rect 554596 702448 554648 702500
rect 559656 702448 559708 702500
rect 8116 700952 8168 701004
rect 13084 700952 13136 701004
rect 40500 700952 40552 701004
rect 44916 700952 44968 701004
rect 56784 700952 56836 701004
rect 60740 700952 60792 701004
rect 72976 700952 73028 701004
rect 76748 700952 76800 701004
rect 89168 700952 89220 701004
rect 92572 700952 92624 701004
rect 105452 700952 105504 701004
rect 108580 700952 108632 701004
rect 121644 700952 121696 701004
rect 124404 700952 124456 701004
rect 137836 700952 137888 701004
rect 140412 700952 140464 701004
rect 154120 700952 154172 701004
rect 156236 700952 156288 701004
rect 170312 700952 170364 701004
rect 172428 700952 172480 701004
rect 202788 700952 202840 701004
rect 204260 700952 204312 701004
rect 348056 700952 348108 701004
rect 348792 700952 348844 701004
rect 363880 700952 363932 701004
rect 364984 700952 365036 701004
rect 379336 700952 379388 701004
rect 381176 700952 381228 701004
rect 395712 700952 395764 701004
rect 397460 700952 397512 701004
rect 411720 700952 411772 701004
rect 413652 700952 413704 701004
rect 427544 700952 427596 701004
rect 429844 700952 429896 701004
rect 443552 700952 443604 701004
rect 446128 700952 446180 701004
rect 475384 700952 475436 701004
rect 478512 700952 478564 701004
rect 59728 3816 59780 3868
rect 74724 3952 74776 4004
rect 58808 3680 58860 3732
rect 70216 3884 70268 3936
rect 62028 3748 62080 3800
rect 67456 3748 67508 3800
rect 78036 3884 78088 3936
rect 63224 3612 63276 3664
rect 69020 3680 69072 3732
rect 71412 3680 71464 3732
rect 69112 3612 69164 3664
rect 83556 3816 83608 3868
rect 80888 3748 80940 3800
rect 94596 3816 94648 3868
rect 122288 3816 122340 3868
rect 133236 3816 133288 3868
rect 84476 3748 84528 3800
rect 98000 3748 98052 3800
rect 114008 3748 114060 3800
rect 125508 3748 125560 3800
rect 66720 3544 66772 3596
rect 81348 3680 81400 3732
rect 85672 3680 85724 3732
rect 56048 3476 56100 3528
rect 69020 3476 69072 3528
rect 70124 3476 70176 3528
rect 54944 3408 54996 3460
rect 70216 3408 70268 3460
rect 72976 3476 73028 3528
rect 86868 3612 86920 3664
rect 87788 3680 87840 3732
rect 101220 3680 101272 3732
rect 116400 3680 116452 3732
rect 127716 3680 127768 3732
rect 99012 3612 99064 3664
rect 109408 3612 109460 3664
rect 121184 3612 121236 3664
rect 125048 3612 125100 3664
rect 135444 3612 135496 3664
rect 143632 3612 143684 3664
rect 153108 3612 153160 3664
rect 82912 3544 82964 3596
rect 83280 3544 83332 3596
rect 96804 3544 96856 3596
rect 102232 3544 102284 3596
rect 114468 3544 114520 3596
rect 121092 3544 121144 3596
rect 132132 3544 132184 3596
rect 136456 3544 136508 3596
rect 146484 3544 146536 3596
rect 149520 3544 149572 3596
rect 158628 3544 158680 3596
rect 78588 3476 78640 3528
rect 92388 3476 92440 3528
rect 51356 3340 51408 3392
rect 66996 3340 67048 3392
rect 67456 3340 67508 3392
rect 76932 3340 76984 3392
rect 65524 3272 65576 3324
rect 50160 3204 50212 3256
rect 65892 3204 65944 3256
rect 71504 3272 71556 3324
rect 85764 3408 85816 3460
rect 90364 3408 90416 3460
rect 103612 3476 103664 3528
rect 110512 3476 110564 3528
rect 122380 3476 122432 3528
rect 127072 3476 127124 3528
rect 137652 3476 137704 3528
rect 139216 3476 139268 3528
rect 148692 3476 148744 3528
rect 153016 3476 153068 3528
rect 160192 3476 160244 3528
rect 79692 3340 79744 3392
rect 83004 3340 83056 3392
rect 89536 3340 89588 3392
rect 102324 3408 102376 3460
rect 105728 3408 105780 3460
rect 117780 3408 117832 3460
rect 131764 3408 131816 3460
rect 142252 3408 142304 3460
rect 142528 3408 142580 3460
rect 151728 3408 151780 3460
rect 155776 3408 155828 3460
rect 96252 3340 96304 3392
rect 109040 3340 109092 3392
rect 112812 3340 112864 3392
rect 124128 3340 124180 3392
rect 125968 3340 126020 3392
rect 136640 3340 136692 3392
rect 82912 3272 82964 3324
rect 84660 3272 84712 3324
rect 86868 3272 86920 3324
rect 100116 3272 100168 3324
rect 103336 3272 103388 3324
rect 115572 3272 115624 3324
rect 117596 3272 117648 3324
rect 128820 3272 128872 3324
rect 129372 3272 129424 3324
rect 139860 3272 139912 3324
rect 149796 3340 149848 3392
rect 148324 3272 148376 3324
rect 157248 3272 157300 3324
rect 79968 3204 80020 3256
rect 93952 3204 94004 3256
rect 106740 3204 106792 3256
rect 107200 3204 107252 3256
rect 118608 3204 118660 3256
rect 119896 3204 119948 3256
rect 131028 3204 131080 3256
rect 140044 3204 140096 3256
rect 154028 3204 154080 3256
rect 40960 3136 41012 3188
rect 57060 3136 57112 3188
rect 57520 3136 57572 3188
rect 72516 3136 72568 3188
rect 73804 3136 73856 3188
rect 87972 3136 88024 3188
rect 101036 3136 101088 3188
rect 113088 3136 113140 3188
rect 52552 3068 52604 3120
rect 68100 3068 68152 3120
rect 76288 3068 76340 3120
rect 44272 3000 44324 3052
rect 60372 3000 60424 3052
rect 64328 3000 64380 3052
rect 79140 3000 79192 3052
rect 79600 3068 79652 3120
rect 89076 3068 89128 3120
rect 98736 3068 98788 3120
rect 111156 3068 111208 3120
rect 111616 3068 111668 3120
rect 123300 3068 123352 3120
rect 33600 2932 33652 2984
rect 50436 2932 50488 2984
rect 26608 2864 26660 2916
rect 43812 2864 43864 2916
rect 48964 2864 49016 2916
rect 64880 2932 64932 2984
rect 67916 2932 67968 2984
rect 82728 2932 82780 2984
rect 83004 3000 83056 3052
rect 93492 3000 93544 3052
rect 95148 3000 95200 3052
rect 107844 3000 107896 3052
rect 108488 3000 108540 3052
rect 119988 3000 120040 3052
rect 134340 3136 134392 3188
rect 137652 3136 137704 3188
rect 147772 3136 147824 3188
rect 134156 3068 134208 3120
rect 144276 3068 144328 3120
rect 147128 3068 147180 3120
rect 156420 3136 156472 3188
rect 128176 3000 128228 3052
rect 138756 3000 138808 3052
rect 90456 2932 90508 2984
rect 91560 2932 91612 2984
rect 104532 2932 104584 2984
rect 104624 2932 104676 2984
rect 116952 2932 117004 2984
rect 123484 2932 123536 2984
rect 130568 2932 130620 2984
rect 140964 2932 141016 2984
rect 27712 2796 27764 2848
rect 45192 2796 45244 2848
rect 47860 2796 47912 2848
rect 63684 2864 63736 2916
rect 75368 2864 75420 2916
rect 79600 2864 79652 2916
rect 82084 2864 82136 2916
rect 95976 2864 96028 2916
rect 97448 2864 97500 2916
rect 110052 2864 110104 2916
rect 115204 2864 115256 2916
rect 126888 2864 126940 2916
rect 132960 2864 133012 2916
rect 143172 3000 143224 3052
rect 145932 3000 145984 3052
rect 155316 3068 155368 3120
rect 166080 3408 166132 3460
rect 158168 3272 158220 3324
rect 166356 3340 166408 3392
rect 174084 3340 174136 3392
rect 161296 3272 161348 3324
rect 169668 3272 169720 3324
rect 181812 3272 181864 3324
rect 564348 3272 564400 3324
rect 583392 3272 583444 3324
rect 160192 3204 160244 3256
rect 161940 3204 161992 3256
rect 163688 3204 163740 3256
rect 171876 3204 171928 3256
rect 174268 3204 174320 3256
rect 164148 3136 164200 3188
rect 170772 3136 170824 3188
rect 178500 3136 178552 3188
rect 162768 3068 162820 3120
rect 164884 3068 164936 3120
rect 172980 3068 173032 3120
rect 173440 3068 173492 3120
rect 180892 3204 180944 3256
rect 184940 3204 184992 3256
rect 181444 3136 181496 3188
rect 188436 3136 188488 3188
rect 200304 3204 200356 3256
rect 206100 3204 206152 3256
rect 556712 3204 556764 3256
rect 575112 3204 575164 3256
rect 191748 3136 191800 3188
rect 195612 3136 195664 3188
rect 201684 3136 201736 3188
rect 220268 3136 220320 3188
rect 224868 3136 224920 3188
rect 561128 3136 561180 3188
rect 579804 3136 579856 3188
rect 179052 3068 179104 3120
rect 186320 3068 186372 3120
rect 190552 3068 190604 3120
rect 197268 3068 197320 3120
rect 202696 3068 202748 3120
rect 208308 3068 208360 3120
rect 209872 3068 209924 3120
rect 214932 3068 214984 3120
rect 215668 3068 215720 3120
rect 220452 3068 220504 3120
rect 221556 3068 221608 3120
rect 225972 3068 226024 3120
rect 228732 3068 228784 3120
rect 232596 3068 232648 3120
rect 239312 3068 239364 3120
rect 242532 3068 242584 3120
rect 543464 3068 543516 3120
rect 560484 3068 560536 3120
rect 562232 3068 562284 3120
rect 581000 3068 581052 3120
rect 151820 3000 151872 3052
rect 160836 3000 160888 3052
rect 162492 3000 162544 3052
rect 170864 3000 170916 3052
rect 171968 3000 172020 3052
rect 179604 3000 179656 3052
rect 182548 3000 182600 3052
rect 189540 3000 189592 3052
rect 189724 3000 189776 3052
rect 196164 3000 196216 3052
rect 141240 2932 141292 2984
rect 150900 2932 150952 2984
rect 156604 2932 156656 2984
rect 165528 2932 165580 2984
rect 167184 2932 167236 2984
rect 175464 2932 175516 2984
rect 175832 2932 175884 2984
rect 144736 2864 144788 2916
rect 60832 2796 60884 2848
rect 75828 2796 75880 2848
rect 77392 2796 77444 2848
rect 91284 2796 91336 2848
rect 92756 2796 92808 2848
rect 98644 2796 98696 2848
rect 99840 2796 99892 2848
rect 112536 2796 112588 2848
rect 118792 2796 118844 2848
rect 130200 2796 130252 2848
rect 135260 2796 135312 2848
rect 145380 2796 145432 2848
rect 150624 2864 150676 2916
rect 160008 2864 160060 2916
rect 160100 2864 160152 2916
rect 168840 2864 168892 2916
rect 169576 2864 169628 2916
rect 177672 2864 177724 2916
rect 177856 2932 177908 2984
rect 185400 2932 185452 2984
rect 194416 2932 194468 2984
rect 200580 3000 200632 3052
rect 203892 3000 203944 3052
rect 209412 3000 209464 3052
rect 212172 3000 212224 3052
rect 217140 3000 217192 3052
rect 219256 3000 219308 3052
rect 223488 3000 223540 3052
rect 228180 3000 228232 3052
rect 229836 3000 229888 3052
rect 233700 3000 233752 3052
rect 234620 3000 234672 3052
rect 238116 3000 238168 3052
rect 240508 3000 240560 3052
rect 243636 3000 243688 3052
rect 245200 3000 245252 3052
rect 248052 3000 248104 3052
rect 248788 3000 248840 3052
rect 251364 3000 251416 3052
rect 333704 3000 333756 3052
rect 336280 3000 336332 3052
rect 530032 3000 530084 3052
rect 546684 3000 546736 3052
rect 553308 3000 553360 3052
rect 571524 3000 571576 3052
rect 199108 2932 199160 2984
rect 204996 2932 205048 2984
rect 182916 2864 182968 2916
rect 183744 2864 183796 2916
rect 190644 2864 190696 2916
rect 192392 2864 192444 2916
rect 198372 2864 198424 2916
rect 201500 2864 201552 2916
rect 206928 2932 206980 2984
rect 208584 2932 208636 2984
rect 213828 2932 213880 2984
rect 214472 2932 214524 2984
rect 219348 2932 219400 2984
rect 223948 2932 224000 2984
rect 225144 2932 225196 2984
rect 229560 2932 229612 2984
rect 231032 2932 231084 2984
rect 235080 2932 235132 2984
rect 235816 2932 235868 2984
rect 239496 2932 239548 2984
rect 242072 2932 242124 2984
rect 245016 2932 245068 2984
rect 247592 2932 247644 2984
rect 250536 2932 250588 2984
rect 253480 2932 253532 2984
rect 256056 2932 256108 2984
rect 310244 2932 310296 2984
rect 311440 2932 311492 2984
rect 325700 2932 325752 2984
rect 328000 2932 328052 2984
rect 329012 2932 329064 2984
rect 331588 2932 331640 2984
rect 332324 2932 332376 2984
rect 335084 2932 335136 2984
rect 341156 2932 341208 2984
rect 344560 2932 344612 2984
rect 513288 2932 513340 2984
rect 529020 2932 529072 2984
rect 549812 2932 549864 2984
rect 568028 2932 568080 2984
rect 206192 2864 206244 2916
rect 211620 2864 211672 2916
rect 213368 2864 213420 2916
rect 217968 2864 218020 2916
rect 218060 2864 218112 2916
rect 222936 2864 222988 2916
rect 223120 2864 223172 2916
rect 227352 2864 227404 2916
rect 227536 2864 227588 2916
rect 231768 2864 231820 2916
rect 232228 2864 232280 2916
rect 236184 2864 236236 2916
rect 237012 2864 237064 2916
rect 240600 2864 240652 2916
rect 244096 2864 244148 2916
rect 247224 2864 247276 2916
rect 249984 2864 250036 2916
rect 252744 2864 252796 2916
rect 254676 2864 254728 2916
rect 257160 2864 257212 2916
rect 261760 2864 261812 2916
rect 263784 2864 263836 2916
rect 312452 2864 312504 2916
rect 313832 2864 313884 2916
rect 314568 2864 314620 2916
rect 316224 2864 316276 2916
rect 316868 2864 316920 2916
rect 318524 2864 318576 2916
rect 319076 2864 319128 2916
rect 320916 2864 320968 2916
rect 321284 2864 321336 2916
rect 323308 2864 323360 2916
rect 323492 2864 323544 2916
rect 325608 2864 325660 2916
rect 327908 2864 327960 2916
rect 330392 2864 330444 2916
rect 331128 2864 331180 2916
rect 333888 2864 333940 2916
rect 334532 2864 334584 2916
rect 337476 2864 337528 2916
rect 340052 2864 340104 2916
rect 342996 2864 343048 2916
rect 517520 2864 517572 2916
rect 523040 2864 523092 2916
rect 525800 2864 525852 2916
rect 531320 2864 531372 2916
rect 536564 2864 536616 2916
rect 553768 2864 553820 2916
rect 559748 2864 559800 2916
rect 578608 2864 578660 2916
rect 154212 2796 154264 2848
rect 158904 2796 158956 2848
rect 167736 2796 167788 2848
rect 168380 2796 168432 2848
rect 176292 2796 176344 2848
rect 180248 2796 180300 2848
rect 187332 2796 187384 2848
rect 199476 2796 199528 2848
rect 205088 2796 205140 2848
rect 210516 2796 210568 2848
rect 210976 2796 211028 2848
rect 216036 2796 216088 2848
rect 216864 2796 216916 2848
rect 221832 2796 221884 2848
rect 226340 2796 226392 2848
rect 230664 2796 230716 2848
rect 233424 2796 233476 2848
rect 237288 2796 237340 2848
rect 238116 2796 238168 2848
rect 241704 2796 241756 2848
rect 242900 2796 242952 2848
rect 246120 2796 246172 2848
rect 246396 2796 246448 2848
rect 249432 2796 249484 2848
rect 252376 2796 252428 2848
rect 254952 2796 255004 2848
rect 255872 2796 255924 2848
rect 258264 2796 258316 2848
rect 260656 2796 260708 2848
rect 262680 2796 262732 2848
rect 304724 2796 304776 2848
rect 305552 2796 305604 2848
rect 306932 2796 306984 2848
rect 307944 2796 307996 2848
rect 309140 2796 309192 2848
rect 310244 2796 310296 2848
rect 311348 2796 311400 2848
rect 312636 2796 312688 2848
rect 313556 2796 313608 2848
rect 315028 2796 315080 2848
rect 315764 2796 315816 2848
rect 317328 2796 317380 2848
rect 317972 2796 318024 2848
rect 319720 2796 319772 2848
rect 320088 2796 320140 2848
rect 322112 2796 322164 2848
rect 322388 2796 322440 2848
rect 324412 2796 324464 2848
rect 324596 2796 324648 2848
rect 326804 2796 326856 2848
rect 326988 2796 327040 2848
rect 329196 2796 329248 2848
rect 330116 2796 330168 2848
rect 332692 2796 332744 2848
rect 335636 2796 335688 2848
rect 338672 2796 338724 2848
rect 338948 2796 339000 2848
rect 342076 2796 342128 2848
rect 346676 2796 346728 2848
rect 350448 2796 350500 2848
rect 353208 2796 353260 2848
rect 357532 2796 357584 2848
rect 372344 2796 372396 2848
rect 377680 2796 377732 2848
rect 517612 2796 517664 2848
rect 521844 2796 521896 2848
rect 562968 2796 563020 2848
rect 582196 2796 582248 2848
rect 193220 2728 193272 2780
rect 176660 1300 176712 1352
rect 184296 1300 184348 1352
rect 187332 1300 187384 1352
rect 194232 1300 194284 1352
rect 198280 1300 198332 1352
rect 204168 1300 204220 1352
rect 207388 1300 207440 1352
rect 213000 1300 213052 1352
rect 257068 1300 257120 1352
rect 259368 1300 259420 1352
rect 259460 1300 259512 1352
rect 261576 1300 261628 1352
rect 262956 1300 263008 1352
rect 264888 1300 264940 1352
rect 265348 1300 265400 1352
rect 267096 1300 267148 1352
rect 267740 1300 267792 1352
rect 269304 1300 269356 1352
rect 271236 1300 271288 1352
rect 272616 1300 272668 1352
rect 273628 1300 273680 1352
rect 274824 1300 274876 1352
rect 277124 1300 277176 1352
rect 278136 1300 278188 1352
rect 279516 1300 279568 1352
rect 280344 1300 280396 1352
rect 336648 1300 336700 1352
rect 339868 1300 339920 1352
rect 342168 1300 342220 1352
rect 345756 1300 345808 1352
rect 348884 1300 348936 1352
rect 352840 1300 352892 1352
rect 356612 1300 356664 1352
rect 361120 1300 361172 1352
rect 364248 1300 364300 1352
rect 369400 1300 369452 1352
rect 374276 1300 374328 1352
rect 379612 1300 379664 1352
rect 384212 1300 384264 1352
rect 390652 1300 390704 1352
rect 396356 1300 396408 1352
rect 403624 1300 403676 1352
rect 406292 1300 406344 1352
rect 414296 1300 414348 1352
rect 419448 1300 419500 1352
rect 428280 1300 428332 1352
rect 428372 1300 428424 1352
rect 98644 1232 98696 1284
rect 105912 1232 105964 1284
rect 188896 1232 188948 1284
rect 195336 1232 195388 1284
rect 197176 1232 197228 1284
rect 203064 1232 203116 1284
rect 258264 1232 258316 1284
rect 260472 1232 260524 1284
rect 264152 1232 264204 1284
rect 265992 1232 266044 1284
rect 266544 1232 266596 1284
rect 268200 1232 268252 1284
rect 270040 1232 270092 1284
rect 271512 1232 271564 1284
rect 272432 1232 272484 1284
rect 273720 1232 273772 1284
rect 343364 1232 343416 1284
rect 346952 1232 347004 1284
rect 349988 1232 350040 1284
rect 354036 1232 354088 1284
rect 357716 1232 357768 1284
rect 362316 1232 362368 1284
rect 365444 1232 365496 1284
rect 370228 1232 370280 1284
rect 370964 1232 371016 1284
rect 376116 1232 376168 1284
rect 377588 1232 377640 1284
rect 383568 1232 383620 1284
rect 388628 1232 388680 1284
rect 395344 1232 395396 1284
rect 404084 1232 404136 1284
rect 411904 1232 411956 1284
rect 413928 1232 413980 1284
rect 422576 1232 422628 1284
rect 426164 1232 426216 1284
rect 435180 1232 435232 1284
rect 436008 1300 436060 1352
rect 437572 1232 437624 1284
rect 438308 1232 438360 1284
rect 443828 1300 443880 1352
rect 454132 1300 454184 1352
rect 186136 1164 186188 1216
rect 193128 1164 193180 1216
rect 268844 1164 268896 1216
rect 270408 1164 270460 1216
rect 359924 1164 359976 1216
rect 364616 1164 364668 1216
rect 366548 1164 366600 1216
rect 371332 1164 371384 1216
rect 378692 1164 378744 1216
rect 384396 1164 384448 1216
rect 387524 1164 387576 1216
rect 394240 1164 394292 1216
rect 395252 1164 395304 1216
rect 402520 1164 402572 1216
rect 412916 1164 412968 1216
rect 421380 1164 421432 1216
rect 421748 1164 421800 1216
rect 430856 1164 430908 1216
rect 439412 1164 439464 1216
rect 443552 1164 443604 1216
rect 445852 1232 445904 1284
rect 449348 1232 449400 1284
rect 456984 1300 457036 1352
rect 457076 1300 457128 1352
rect 468300 1300 468352 1352
rect 481364 1300 481416 1352
rect 494704 1300 494756 1352
rect 495716 1300 495768 1352
rect 509700 1300 509752 1352
rect 510068 1300 510120 1352
rect 525432 1300 525484 1352
rect 539876 1300 539928 1352
rect 556988 1300 557040 1352
rect 454868 1232 454920 1284
rect 448612 1164 448664 1216
rect 450452 1164 450504 1216
rect 462596 1232 462648 1284
rect 474188 1232 474240 1284
rect 480168 1232 480220 1284
rect 493140 1232 493192 1284
rect 493508 1232 493560 1284
rect 507308 1232 507360 1284
rect 507768 1232 507820 1284
rect 517520 1232 517572 1284
rect 534356 1232 534408 1284
rect 551100 1232 551152 1284
rect 352196 1096 352248 1148
rect 356336 1096 356388 1148
rect 361028 1096 361080 1148
rect 365444 1096 365496 1148
rect 367652 1096 367704 1148
rect 372896 1096 372948 1148
rect 375288 1096 375340 1148
rect 4068 1028 4120 1080
rect 23112 1028 23164 1080
rect 355508 1028 355560 1080
rect 359924 1028 359976 1080
rect 373172 1028 373224 1080
rect 378508 1028 378560 1080
rect 379796 1096 379848 1148
rect 385960 1096 386012 1148
rect 386328 1096 386380 1148
rect 392676 1096 392728 1148
rect 397368 1096 397420 1148
rect 404820 1096 404872 1148
rect 420644 1096 420696 1148
rect 429292 1096 429344 1148
rect 434996 1096 435048 1148
rect 445024 1096 445076 1148
rect 445208 1096 445260 1148
rect 455696 1096 455748 1148
rect 465908 1164 465960 1216
rect 475844 1164 475896 1216
rect 488816 1164 488868 1216
rect 501236 1164 501288 1216
rect 515496 1164 515548 1216
rect 516692 1164 516744 1216
rect 532056 1164 532108 1216
rect 461584 1096 461636 1148
rect 469128 1096 469180 1148
rect 481364 1096 481416 1148
rect 487988 1096 488040 1148
rect 501420 1096 501472 1148
rect 506756 1096 506808 1148
rect 517612 1096 517664 1148
rect 522212 1096 522264 1148
rect 538128 1096 538180 1148
rect 381176 1028 381228 1080
rect 385316 1028 385368 1080
rect 391848 1028 391900 1080
rect 394148 1028 394200 1080
rect 401324 1028 401376 1080
rect 415124 1028 415176 1080
rect 423404 1028 423456 1080
rect 424968 1028 425020 1080
rect 434076 1028 434128 1080
rect 441528 1028 441580 1080
rect 451740 1028 451792 1080
rect 455972 1028 456024 1080
rect 467472 1028 467524 1080
rect 474648 1028 474700 1080
rect 487252 1028 487304 1080
rect 518808 1028 518860 1080
rect 534540 1028 534592 1080
rect 20628 960 20680 1012
rect 38568 960 38620 1012
rect 345572 960 345624 1012
rect 349252 960 349304 1012
rect 351092 960 351144 1012
rect 355232 960 355284 1012
rect 362132 960 362184 1012
rect 367008 960 367060 1012
rect 369768 960 369820 1012
rect 375288 960 375340 1012
rect 376484 960 376536 1012
rect 382372 960 382424 1012
rect 422852 960 422904 1012
rect 431868 960 431920 1012
rect 432788 960 432840 1012
rect 442632 960 442684 1012
rect 443552 960 443604 1012
rect 449808 960 449860 1012
rect 489092 960 489144 1012
rect 502984 960 503036 1012
rect 520004 960 520056 1012
rect 536104 960 536156 1012
rect 1676 892 1728 944
rect 20904 892 20956 944
rect 358728 892 358780 944
rect 363512 892 363564 944
rect 416228 892 416280 944
rect 424968 892 425020 944
rect 433892 892 433944 944
rect 443460 892 443512 944
rect 446036 892 446088 944
rect 456892 892 456944 944
rect 494612 892 494664 944
rect 508872 892 508924 944
rect 515588 892 515640 944
rect 525800 892 525852 944
rect 532148 892 532200 944
rect 548708 892 548760 944
rect 19432 824 19484 876
rect 37464 824 37516 876
rect 337844 824 337896 876
rect 340972 824 341024 876
rect 347688 824 347740 876
rect 351644 824 351696 876
rect 368756 824 368808 876
rect 373908 824 373960 876
rect 448244 824 448296 876
rect 459192 824 459244 876
rect 485688 824 485740 876
rect 498936 824 498988 876
rect 527732 824 527784 876
rect 544384 824 544436 876
rect 547604 824 547656 876
rect 565636 824 565688 876
rect 18236 756 18288 808
rect 36360 756 36412 808
rect 251180 756 251232 808
rect 253848 756 253900 808
rect 427268 756 427320 808
rect 436744 756 436796 808
rect 442724 756 442776 808
rect 453304 756 453356 808
rect 9956 688 10008 740
rect 28632 688 28684 740
rect 401876 688 401928 740
rect 409236 688 409288 740
rect 429476 688 429528 740
rect 439136 688 439188 740
rect 440516 688 440568 740
rect 450912 688 450964 740
rect 451556 688 451608 740
rect 462412 756 462464 808
rect 483572 756 483624 808
rect 497096 756 497148 808
rect 499028 756 499080 808
rect 513564 756 513616 808
rect 528836 756 528888 808
rect 545488 756 545540 808
rect 550916 756 550968 808
rect 569132 756 569184 808
rect 468116 688 468168 740
rect 480536 688 480588 740
rect 482468 688 482520 740
rect 495532 688 495584 740
rect 502248 688 502300 740
rect 517152 688 517204 740
rect 521108 688 521160 740
rect 537208 688 537260 740
rect 537668 688 537720 740
rect 554964 688 555016 740
rect 8760 620 8812 672
rect 27528 620 27580 672
rect 34796 620 34848 672
rect 51816 620 51868 672
rect 393044 620 393096 672
rect 400128 620 400180 672
rect 400772 620 400824 672
rect 408592 620 408644 672
rect 409604 620 409656 672
rect 417884 620 417936 672
rect 14740 552 14792 604
rect 17040 552 17092 604
rect 35256 552 35308 604
rect 35992 552 36044 604
rect 52920 552 52972 604
rect 389732 552 389784 604
rect 396540 552 396592 604
rect 408408 552 408460 604
rect 416688 552 416740 604
rect 431684 552 431736 604
rect 441528 620 441580 672
rect 456984 620 457036 672
rect 460020 620 460072 672
rect 464804 620 464856 672
rect 476948 620 477000 672
rect 486884 620 486936 672
rect 500592 620 500644 672
rect 503444 620 503496 672
rect 518348 620 518400 672
rect 523316 620 523368 672
rect 33048 484 33100 536
rect 39764 484 39816 536
rect 56232 484 56284 536
rect 430488 484 430540 536
rect 440332 552 440384 604
rect 447048 552 447100 604
rect 458088 552 458140 604
rect 461492 552 461544 604
rect 473452 552 473504 604
rect 486424 552 486476 604
rect 459468 484 459520 536
rect 470784 484 470836 536
rect 473636 484 473688 536
rect 16212 416 16264 468
rect 34152 416 34204 468
rect 38568 416 38620 468
rect 55128 416 55180 468
rect 382004 416 382056 468
rect 387892 416 387944 468
rect 412088 416 412140 468
rect 420368 416 420420 468
rect 437204 416 437256 468
rect 447232 416 447284 468
rect 470324 416 470376 468
rect 482468 416 482520 468
rect 484676 416 484728 468
rect 498200 552 498252 604
rect 490196 416 490248 468
rect 503812 552 503864 604
rect 508964 552 509016 604
rect 523868 552 523920 604
rect 524328 620 524380 672
rect 533252 620 533304 672
rect 539600 620 539652 672
rect 542084 620 542136 672
rect 533712 552 533764 604
rect 533804 552 533856 604
rect 11520 348 11572 400
rect 29736 348 29788 400
rect 32220 348 32272 400
rect 49608 348 49660 400
rect 407396 348 407448 400
rect 415308 348 415360 400
rect 460572 348 460624 400
rect 472440 348 472492 400
rect 478328 348 478380 400
rect 490748 348 490800 400
rect 497924 348 497976 400
rect 512092 484 512144 536
rect 517796 484 517848 536
rect 500132 416 500184 468
rect 514944 416 514996 468
rect 525708 416 525760 468
rect 542176 416 542228 468
rect 504548 348 504600 400
rect 519728 348 519780 400
rect 533252 348 533304 400
rect 540428 348 540480 400
rect 548984 620 549036 672
rect 566832 620 566884 672
rect 545396 552 545448 604
rect 563244 552 563296 604
rect 559380 484 559432 536
rect 544568 416 544620 468
rect 562232 416 562284 468
rect 550456 348 550508 400
rect 555332 348 555384 400
rect 573548 348 573600 400
rect 3240 280 3292 332
rect 22008 280 22060 332
rect 30288 280 30340 332
rect 47400 280 47452 332
rect 398564 280 398616 332
rect 406200 280 406252 332
rect 410984 280 411036 332
rect 418620 280 418672 332
rect 453764 280 453816 332
rect 464988 280 465040 332
rect 471428 280 471480 332
rect 484216 280 484268 332
rect 505652 280 505704 332
rect 520372 280 520424 332
rect 531044 280 531096 332
rect 548064 280 548116 332
rect 551928 280 551980 332
rect 570512 280 570564 332
rect 22836 212 22888 264
rect 40500 212 40552 264
rect 42248 212 42300 264
rect 58164 212 58216 264
rect 354404 212 354456 264
rect 358912 212 358964 264
rect 380808 212 380860 264
rect 386788 212 386840 264
rect 391664 212 391716 264
rect 398748 212 398800 264
rect 405188 212 405240 264
rect 412824 212 412876 264
rect 457904 212 457956 264
rect 470048 212 470100 264
rect 472532 212 472584 264
rect 484860 212 484912 264
rect 511448 212 511500 264
rect 526260 212 526312 264
rect 538772 212 538824 264
rect 556344 212 556396 264
rect 557172 212 557224 264
rect 575940 212 575992 264
rect 8024 144 8076 196
rect 26332 144 26384 196
rect 31116 144 31168 196
rect 48504 144 48556 196
rect 53564 144 53616 196
rect 69480 144 69532 196
rect 418436 144 418488 196
rect 426900 144 426952 196
rect 465816 144 465868 196
rect 478328 144 478380 196
rect 479156 144 479208 196
rect 492496 144 492548 196
rect 492588 144 492640 196
rect 506664 144 506716 196
rect 512644 144 512696 196
rect 528008 144 528060 196
rect 535368 144 535420 196
rect 552848 144 552900 196
rect 554228 144 554280 196
rect 572904 144 572956 196
rect 22008 76 22060 128
rect 39396 76 39448 128
rect 45284 76 45336 128
rect 61752 76 61804 128
rect 399668 76 399720 128
rect 407028 76 407080 128
rect 423956 76 424008 128
rect 433432 76 433484 128
rect 452568 76 452620 128
rect 464160 76 464212 128
rect 467012 76 467064 128
rect 478972 76 479024 128
rect 491300 76 491352 128
rect 505560 76 505612 128
rect 514484 76 514536 128
rect 529940 76 529992 128
rect 540980 76 541032 128
rect 558736 76 558788 128
rect 558828 76 558880 128
rect 577136 76 577188 128
rect 388 8 440 60
rect 19800 8 19852 60
rect 24584 8 24636 60
rect 41604 8 41656 60
rect 42892 8 42944 60
rect 59360 8 59412 60
rect 344744 8 344796 60
rect 348240 8 348292 60
rect 363236 8 363288 60
rect 367836 8 367888 60
rect 383108 8 383160 60
rect 389640 8 389692 60
rect 390836 8 390888 60
rect 397920 8 397972 60
rect 402888 8 402940 60
rect 410984 8 411036 60
rect 417332 8 417384 60
rect 425796 8 425848 60
rect 463608 8 463660 60
rect 475936 8 475988 60
rect 477224 8 477276 60
rect 490104 8 490156 60
rect 496728 8 496780 60
rect 511448 8 511500 60
rect 526904 8 526956 60
rect 542820 8 542872 60
rect 546408 8 546460 60
rect 564624 8 564676 60
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 251652 703582 251864 703610
rect 8128 701010 8156 703520
rect 24320 702506 24348 703520
rect 24308 702500 24360 702506
rect 24308 702442 24360 702448
rect 29276 702500 29328 702506
rect 29276 702442 29328 702448
rect 8116 701004 8168 701010
rect 8116 700946 8168 700952
rect 13084 701004 13136 701010
rect 13084 700946 13136 700952
rect 13096 700890 13124 700946
rect 13096 700862 13386 700890
rect 29288 700876 29316 702442
rect 40512 701010 40540 703520
rect 56796 701010 56824 703520
rect 72988 701010 73016 703520
rect 89180 701010 89208 703520
rect 105464 701010 105492 703520
rect 121656 701010 121684 703520
rect 137848 701010 137876 703520
rect 154132 701010 154160 703520
rect 170324 701010 170352 703520
rect 186516 703050 186544 703520
rect 186504 703044 186556 703050
rect 186504 702986 186556 702992
rect 188436 703044 188488 703050
rect 188436 702986 188488 702992
rect 40500 701004 40552 701010
rect 40500 700946 40552 700952
rect 44916 701004 44968 701010
rect 44916 700946 44968 700952
rect 56784 701004 56836 701010
rect 56784 700946 56836 700952
rect 60740 701004 60792 701010
rect 60740 700946 60792 700952
rect 72976 701004 73028 701010
rect 72976 700946 73028 700952
rect 76748 701004 76800 701010
rect 76748 700946 76800 700952
rect 89168 701004 89220 701010
rect 89168 700946 89220 700952
rect 92572 701004 92624 701010
rect 92572 700946 92624 700952
rect 105452 701004 105504 701010
rect 105452 700946 105504 700952
rect 108580 701004 108632 701010
rect 108580 700946 108632 700952
rect 121644 701004 121696 701010
rect 121644 700946 121696 700952
rect 124404 701004 124456 701010
rect 124404 700946 124456 700952
rect 137836 701004 137888 701010
rect 137836 700946 137888 700952
rect 140412 701004 140464 701010
rect 140412 700946 140464 700952
rect 154120 701004 154172 701010
rect 154120 700946 154172 700952
rect 156236 701004 156288 701010
rect 156236 700946 156288 700952
rect 170312 701004 170364 701010
rect 170312 700946 170364 700952
rect 172428 701004 172480 701010
rect 172428 700946 172480 700952
rect 44928 700890 44956 700946
rect 60752 700890 60780 700946
rect 76760 700890 76788 700946
rect 92584 700890 92612 700946
rect 108592 700890 108620 700946
rect 124416 700890 124444 700946
rect 140424 700890 140452 700946
rect 156248 700890 156276 700946
rect 172440 700890 172468 700946
rect 44928 700862 45218 700890
rect 60752 700862 61134 700890
rect 76760 700862 77050 700890
rect 92584 700862 92966 700890
rect 108592 700862 108882 700890
rect 124416 700862 124798 700890
rect 140424 700862 140714 700890
rect 156248 700862 156630 700890
rect 172440 700862 172546 700890
rect 188448 700876 188476 702986
rect 202800 701010 202828 703520
rect 218992 702506 219020 703520
rect 235184 703050 235212 703520
rect 251468 703474 251496 703520
rect 251652 703474 251680 703582
rect 251468 703446 251680 703474
rect 235172 703044 235224 703050
rect 235172 702986 235224 702992
rect 236184 703044 236236 703050
rect 236184 702986 236236 702992
rect 218980 702500 219032 702506
rect 218980 702442 219032 702448
rect 220268 702500 220320 702506
rect 220268 702442 220320 702448
rect 202788 701004 202840 701010
rect 202788 700946 202840 700952
rect 204260 701004 204312 701010
rect 204260 700946 204312 700952
rect 204272 700890 204300 700946
rect 204272 700862 204378 700890
rect 220280 700876 220308 702442
rect 236196 700876 236224 702986
rect 251836 700890 251864 703582
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332152 703582 332364 703610
rect 267660 700890 267688 703520
rect 283852 700890 283880 703520
rect 300136 700890 300164 703520
rect 316328 702434 316356 703520
rect 316052 702406 316356 702434
rect 316052 700890 316080 702406
rect 332152 700890 332180 703582
rect 332336 703474 332364 703582
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 332520 703474 332548 703520
rect 332336 703446 332548 703474
rect 348804 701010 348832 703520
rect 364996 701010 365024 703520
rect 381188 701010 381216 703520
rect 397472 701010 397500 703520
rect 413664 701010 413692 703520
rect 429856 701010 429884 703520
rect 446140 701010 446168 703520
rect 462332 702506 462360 703520
rect 459100 702500 459152 702506
rect 459100 702442 459152 702448
rect 462320 702500 462372 702506
rect 462320 702442 462372 702448
rect 348056 701004 348108 701010
rect 348056 700946 348108 700952
rect 348792 701004 348844 701010
rect 348792 700946 348844 700952
rect 363880 701004 363932 701010
rect 363880 700946 363932 700952
rect 364984 701004 365036 701010
rect 364984 700946 365036 700952
rect 379336 701004 379388 701010
rect 379336 700946 379388 700952
rect 381176 701004 381228 701010
rect 381176 700946 381228 700952
rect 395712 701004 395764 701010
rect 395712 700946 395764 700952
rect 397460 701004 397512 701010
rect 397460 700946 397512 700952
rect 411720 701004 411772 701010
rect 411720 700946 411772 700952
rect 413652 701004 413704 701010
rect 413652 700946 413704 700952
rect 427544 701004 427596 701010
rect 427544 700946 427596 700952
rect 429844 701004 429896 701010
rect 429844 700946 429896 700952
rect 443552 701004 443604 701010
rect 443552 700946 443604 700952
rect 446128 701004 446180 701010
rect 446128 700946 446180 700952
rect 348068 700890 348096 700946
rect 363892 700890 363920 700946
rect 251836 700862 252126 700890
rect 267660 700862 268042 700890
rect 283852 700862 283958 700890
rect 299966 700862 300164 700890
rect 315882 700862 316080 700890
rect 331798 700862 332180 700890
rect 347714 700862 348096 700890
rect 363630 700862 363920 700890
rect 379348 700890 379376 700946
rect 395724 700890 395752 700946
rect 411732 700890 411760 700946
rect 427556 700890 427584 700946
rect 443564 700890 443592 700946
rect 379348 700862 379454 700890
rect 395462 700862 395752 700890
rect 411378 700862 411760 700890
rect 427294 700862 427584 700890
rect 443210 700862 443592 700890
rect 459112 700876 459140 702442
rect 478524 701010 478552 703520
rect 494808 702778 494836 703520
rect 490932 702772 490984 702778
rect 490932 702714 490984 702720
rect 494796 702772 494848 702778
rect 494796 702714 494848 702720
rect 475384 701004 475436 701010
rect 475384 700946 475436 700952
rect 478512 701004 478564 701010
rect 478512 700946 478564 700952
rect 475396 700890 475424 700946
rect 475042 700862 475424 700890
rect 490944 700876 490972 702714
rect 511000 702506 511028 703520
rect 527192 703066 527220 703520
rect 527100 703050 527220 703066
rect 522764 703044 522816 703050
rect 522764 702986 522816 702992
rect 527088 703044 527220 703050
rect 527140 703038 527220 703044
rect 527088 702986 527140 702992
rect 506848 702500 506900 702506
rect 506848 702442 506900 702448
rect 510988 702500 511040 702506
rect 510988 702442 511040 702448
rect 506860 700876 506888 702442
rect 522776 700876 522804 702986
rect 543476 702778 543504 703520
rect 538680 702772 538732 702778
rect 538680 702714 538732 702720
rect 543464 702772 543516 702778
rect 543464 702714 543516 702720
rect 538692 700876 538720 702714
rect 559668 702506 559696 703520
rect 575860 703050 575888 703520
rect 570512 703044 570564 703050
rect 570512 702986 570564 702992
rect 575848 703044 575900 703050
rect 575848 702986 575900 702992
rect 554596 702500 554648 702506
rect 554596 702442 554648 702448
rect 559656 702500 559708 702506
rect 559656 702442 559708 702448
rect 554608 700876 554636 702442
rect 570524 700876 570552 702986
rect 2778 697368 2834 697377
rect 2778 697303 2834 697312
rect 2792 690849 2820 697303
rect 581642 697232 581698 697241
rect 581642 697167 581698 697176
rect 581656 691529 581684 697167
rect 581642 691520 581698 691529
rect 581642 691455 581698 691464
rect 2778 690840 2834 690849
rect 2778 690775 2834 690784
rect 2778 684312 2834 684321
rect 2778 684247 2834 684256
rect 2792 678065 2820 684247
rect 582378 683904 582434 683913
rect 582378 683839 582434 683848
rect 582392 678473 582420 683839
rect 582378 678464 582434 678473
rect 582378 678399 582434 678408
rect 2778 678056 2834 678065
rect 2778 677991 2834 678000
rect 2778 671256 2834 671265
rect 2778 671191 2834 671200
rect 2792 665281 2820 671191
rect 582378 670712 582434 670721
rect 582378 670647 582434 670656
rect 582392 665417 582420 670647
rect 582378 665408 582434 665417
rect 582378 665343 582434 665352
rect 2778 665272 2834 665281
rect 2778 665207 2834 665216
rect 2778 658200 2834 658209
rect 2778 658135 2834 658144
rect 2792 652497 2820 658135
rect 582378 657384 582434 657393
rect 582378 657319 582434 657328
rect 2778 652488 2834 652497
rect 2778 652423 2834 652432
rect 582392 652361 582420 657319
rect 582378 652352 582434 652361
rect 582378 652287 582434 652296
rect 2778 645144 2834 645153
rect 2778 645079 2834 645088
rect 2792 639713 2820 645079
rect 581642 644056 581698 644065
rect 581642 643991 581698 644000
rect 2778 639704 2834 639713
rect 2778 639639 2834 639648
rect 581656 639305 581684 643991
rect 581642 639296 581698 639305
rect 581642 639231 581698 639240
rect 2778 632088 2834 632097
rect 2778 632023 2834 632032
rect 2792 626929 2820 632023
rect 582378 630864 582434 630873
rect 582378 630799 582434 630808
rect 2778 626920 2834 626929
rect 2778 626855 2834 626864
rect 582392 626249 582420 630799
rect 582378 626240 582434 626249
rect 582378 626175 582434 626184
rect 2778 619168 2834 619177
rect 2778 619103 2834 619112
rect 2792 614009 2820 619103
rect 581642 617536 581698 617545
rect 581642 617471 581698 617480
rect 2778 614000 2834 614009
rect 2778 613935 2834 613944
rect 581656 613193 581684 617471
rect 581642 613184 581698 613193
rect 581642 613119 581698 613128
rect 2778 606112 2834 606121
rect 2778 606047 2834 606056
rect 2792 601361 2820 606047
rect 581642 604208 581698 604217
rect 581642 604143 581698 604152
rect 2778 601352 2834 601361
rect 2778 601287 2834 601296
rect 581656 600137 581684 604143
rect 581642 600128 581698 600137
rect 581642 600063 581698 600072
rect 1582 593056 1638 593065
rect 1582 592991 1638 593000
rect 1596 588577 1624 592991
rect 581642 591016 581698 591025
rect 581642 590951 581698 590960
rect 1582 588568 1638 588577
rect 1582 588503 1638 588512
rect 581656 587081 581684 590951
rect 581642 587072 581698 587081
rect 581642 587007 581698 587016
rect 2042 580000 2098 580009
rect 2042 579935 2098 579944
rect 2056 575793 2084 579935
rect 581642 577688 581698 577697
rect 581642 577623 581698 577632
rect 2042 575784 2098 575793
rect 2042 575719 2098 575728
rect 581656 574025 581684 577623
rect 581642 574016 581698 574025
rect 581642 573951 581698 573960
rect 1490 566944 1546 566953
rect 1490 566879 1546 566888
rect 1504 563009 1532 566879
rect 582378 564360 582434 564369
rect 582378 564295 582434 564304
rect 1490 563000 1546 563009
rect 1490 562935 1546 562944
rect 582392 560969 582420 564295
rect 582378 560960 582434 560969
rect 582378 560895 582434 560904
rect 1490 553888 1546 553897
rect 1490 553823 1546 553832
rect 1504 550225 1532 553823
rect 581642 551168 581698 551177
rect 581642 551103 581698 551112
rect 1490 550216 1546 550225
rect 1490 550151 1546 550160
rect 581656 547777 581684 551103
rect 581642 547768 581698 547777
rect 581642 547703 581698 547712
rect 1398 540832 1454 540841
rect 1398 540767 1454 540776
rect 1412 537441 1440 540767
rect 582378 537840 582434 537849
rect 582378 537775 582434 537784
rect 1398 537432 1454 537441
rect 1398 537367 1454 537376
rect 582392 534857 582420 537775
rect 582378 534848 582434 534857
rect 582378 534783 582434 534792
rect 1490 527912 1546 527921
rect 1490 527847 1546 527856
rect 1504 524657 1532 527847
rect 1490 524648 1546 524657
rect 1490 524583 1546 524592
rect 582378 524512 582434 524521
rect 582378 524447 582434 524456
rect 582392 521801 582420 524447
rect 582378 521792 582434 521801
rect 582378 521727 582434 521736
rect 1582 514856 1638 514865
rect 1582 514791 1638 514800
rect 1596 511873 1624 514791
rect 1582 511864 1638 511873
rect 1582 511799 1638 511808
rect 582378 511320 582434 511329
rect 582378 511255 582434 511264
rect 582392 508745 582420 511255
rect 582378 508736 582434 508745
rect 582378 508671 582434 508680
rect 1582 501800 1638 501809
rect 1582 501735 1638 501744
rect 1596 499089 1624 501735
rect 1582 499080 1638 499089
rect 1582 499015 1638 499024
rect 581642 497992 581698 498001
rect 581642 497927 581698 497936
rect 581656 495689 581684 497927
rect 581642 495680 581698 495689
rect 581642 495615 581698 495624
rect 1582 488744 1638 488753
rect 1582 488679 1638 488688
rect 1596 486305 1624 488679
rect 1582 486296 1638 486305
rect 1582 486231 1638 486240
rect 582378 484664 582434 484673
rect 582378 484599 582434 484608
rect 582392 482633 582420 484599
rect 582378 482624 582434 482633
rect 582378 482559 582434 482568
rect 2778 475688 2834 475697
rect 2778 475623 2834 475632
rect 2792 473521 2820 475623
rect 2778 473512 2834 473521
rect 2778 473447 2834 473456
rect 581642 471472 581698 471481
rect 581642 471407 581698 471416
rect 581656 469577 581684 471407
rect 581642 469568 581698 469577
rect 581642 469503 581698 469512
rect 1582 462632 1638 462641
rect 1582 462567 1638 462576
rect 1596 460737 1624 462567
rect 1582 460728 1638 460737
rect 1582 460663 1638 460672
rect 581642 458144 581698 458153
rect 581642 458079 581698 458088
rect 581656 456521 581684 458079
rect 581642 456512 581698 456521
rect 581642 456447 581698 456456
rect 2778 449576 2834 449585
rect 2778 449511 2834 449520
rect 2792 447953 2820 449511
rect 2778 447944 2834 447953
rect 2778 447879 2834 447888
rect 2778 436656 2834 436665
rect 2778 436591 2834 436600
rect 2792 435169 2820 436591
rect 2778 435160 2834 435169
rect 2778 435095 2834 435104
rect 2778 423600 2834 423609
rect 2778 423535 2834 423544
rect 2792 422385 2820 423535
rect 2778 422376 2834 422385
rect 2778 422311 2834 422320
rect 1306 294400 1362 294409
rect 1306 294335 1362 294344
rect 1320 293185 1348 294335
rect 1306 293176 1362 293185
rect 1306 293111 1362 293120
rect 2778 281616 2834 281625
rect 2778 281551 2834 281560
rect 2792 280129 2820 281551
rect 2778 280120 2834 280129
rect 2778 280055 2834 280064
rect 1306 268832 1362 268841
rect 1306 268767 1362 268776
rect 1320 267209 1348 268767
rect 1306 267200 1362 267209
rect 1306 267135 1362 267144
rect 582378 260536 582434 260545
rect 582378 260471 582434 260480
rect 582392 258913 582420 260471
rect 582378 258904 582434 258913
rect 582378 258839 582434 258848
rect 1306 256048 1362 256057
rect 1306 255983 1362 255992
rect 1320 254153 1348 255983
rect 1306 254144 1362 254153
rect 1306 254079 1362 254088
rect 580906 247072 580962 247081
rect 580906 247007 580962 247016
rect 580920 245585 580948 247007
rect 580906 245576 580962 245585
rect 580906 245511 580962 245520
rect 2778 243264 2834 243273
rect 2778 243199 2834 243208
rect 2792 241097 2820 243199
rect 2778 241088 2834 241097
rect 2778 241023 2834 241032
rect 582378 234424 582434 234433
rect 582378 234359 582434 234368
rect 582392 232393 582420 234359
rect 582378 232384 582434 232393
rect 582378 232319 582434 232328
rect 2778 230616 2834 230625
rect 2778 230551 2834 230560
rect 2792 228041 2820 230551
rect 2778 228032 2834 228041
rect 2778 227967 2834 227976
rect 580906 220960 580962 220969
rect 580906 220895 580962 220904
rect 580920 219065 580948 220895
rect 580906 219056 580962 219065
rect 580906 218991 580962 219000
rect 2778 217696 2834 217705
rect 2778 217631 2834 217640
rect 2792 214985 2820 217631
rect 2778 214976 2834 214985
rect 2778 214911 2834 214920
rect 582378 208312 582434 208321
rect 582378 208247 582434 208256
rect 582392 205737 582420 208247
rect 582378 205728 582434 205737
rect 582378 205663 582434 205672
rect 2778 204912 2834 204921
rect 2778 204847 2834 204856
rect 2792 201929 2820 204847
rect 2778 201920 2834 201929
rect 2778 201855 2834 201864
rect 580906 194712 580962 194721
rect 580906 194647 580962 194656
rect 580920 192545 580948 194647
rect 580906 192536 580962 192545
rect 580906 192471 580962 192480
rect 1306 192128 1362 192137
rect 1306 192063 1362 192072
rect 1320 188873 1348 192063
rect 1306 188864 1362 188873
rect 1306 188799 1362 188808
rect 580906 182472 580962 182481
rect 580906 182407 580962 182416
rect 2778 179344 2834 179353
rect 2778 179279 2834 179288
rect 2792 175953 2820 179279
rect 580920 179217 580948 182407
rect 580906 179208 580962 179217
rect 580906 179143 580962 179152
rect 2778 175944 2834 175953
rect 2778 175879 2834 175888
rect 580906 168600 580962 168609
rect 580906 168535 580962 168544
rect 2778 166560 2834 166569
rect 2778 166495 2834 166504
rect 2792 162897 2820 166495
rect 580920 165889 580948 168535
rect 580906 165880 580962 165889
rect 580906 165815 580962 165824
rect 2778 162888 2834 162897
rect 2778 162823 2834 162832
rect 580906 156360 580962 156369
rect 580906 156295 580962 156304
rect 1306 153776 1362 153785
rect 1306 153711 1362 153720
rect 1320 149841 1348 153711
rect 580920 152697 580948 156295
rect 580906 152688 580962 152697
rect 580906 152623 580962 152632
rect 1306 149832 1362 149841
rect 1306 149767 1362 149776
rect 580906 142624 580962 142633
rect 580906 142559 580962 142568
rect 570 140992 626 141001
rect 570 140927 626 140936
rect 584 136785 612 140927
rect 580920 139369 580948 142559
rect 580906 139360 580962 139369
rect 580906 139295 580962 139304
rect 570 136776 626 136785
rect 570 136711 626 136720
rect 580906 130248 580962 130257
rect 580906 130183 580962 130192
rect 754 128208 810 128217
rect 754 128143 810 128152
rect 768 123729 796 128143
rect 580920 126041 580948 130183
rect 580906 126032 580962 126041
rect 580906 125967 580962 125976
rect 754 123720 810 123729
rect 754 123655 810 123664
rect 579894 116376 579950 116385
rect 579894 116311 579950 116320
rect 1306 115424 1362 115433
rect 1306 115359 1362 115368
rect 1320 110673 1348 115359
rect 579908 112849 579936 116311
rect 579894 112840 579950 112849
rect 579894 112775 579950 112784
rect 1306 110664 1362 110673
rect 1306 110599 1362 110608
rect 580906 103592 580962 103601
rect 580906 103527 580962 103536
rect 1582 102640 1638 102649
rect 1582 102575 1638 102584
rect 1596 97617 1624 102575
rect 580920 99521 580948 103527
rect 580906 99512 580962 99521
rect 580906 99447 580962 99456
rect 1582 97608 1638 97617
rect 1582 97543 1638 97552
rect 580906 90264 580962 90273
rect 580906 90199 580962 90208
rect 1582 89856 1638 89865
rect 1582 89791 1638 89800
rect 1596 84697 1624 89791
rect 580920 86193 580948 90199
rect 580906 86184 580962 86193
rect 580906 86119 580962 86128
rect 1582 84688 1638 84697
rect 1582 84623 1638 84632
rect 579894 77344 579950 77353
rect 579894 77279 579950 77288
rect 1582 77072 1638 77081
rect 1582 77007 1638 77016
rect 1596 71641 1624 77007
rect 579908 73001 579936 77279
rect 579894 72992 579950 73001
rect 579894 72927 579950 72936
rect 1582 71632 1638 71641
rect 1582 71567 1638 71576
rect 1490 64288 1546 64297
rect 1490 64223 1546 64232
rect 1504 58585 1532 64223
rect 580906 64152 580962 64161
rect 580906 64087 580962 64096
rect 580920 59673 580948 64087
rect 580906 59664 580962 59673
rect 580906 59599 580962 59608
rect 1490 58576 1546 58585
rect 1490 58511 1546 58520
rect 2042 51504 2098 51513
rect 2042 51439 2098 51448
rect 2056 45529 2084 51439
rect 580906 51096 580962 51105
rect 580906 51031 580962 51040
rect 580920 46345 580948 51031
rect 580906 46336 580962 46345
rect 580906 46271 580962 46280
rect 2042 45520 2098 45529
rect 2042 45455 2098 45464
rect 2042 38720 2098 38729
rect 2042 38655 2098 38664
rect 2056 32473 2084 38655
rect 580906 38040 580962 38049
rect 580906 37975 580962 37984
rect 580920 33153 580948 37975
rect 580906 33144 580962 33153
rect 580906 33079 580962 33088
rect 2042 32464 2098 32473
rect 2042 32399 2098 32408
rect 1490 25936 1546 25945
rect 1490 25871 1546 25880
rect 1504 19417 1532 25871
rect 580906 24984 580962 24993
rect 580906 24919 580962 24928
rect 580920 19825 580948 24919
rect 580906 19816 580962 19825
rect 580906 19751 580962 19760
rect 1490 19408 1546 19417
rect 1490 19343 1546 19352
rect 2042 13152 2098 13161
rect 2042 13087 2098 13096
rect 2056 6497 2084 13087
rect 579894 12744 579950 12753
rect 579894 12679 579950 12688
rect 579908 6633 579936 12679
rect 579894 6624 579950 6633
rect 579894 6559 579950 6568
rect 2042 6488 2098 6497
rect 2042 6423 2098 6432
rect 74736 4010 75026 4026
rect 74724 4004 75026 4010
rect 74776 3998 75026 4004
rect 74724 3946 74776 3952
rect 70216 3936 70268 3942
rect 70214 3904 70216 3913
rect 78036 3936 78088 3942
rect 70268 3904 70270 3913
rect 59728 3868 59780 3874
rect 70214 3839 70270 3848
rect 73618 3904 73674 3913
rect 73674 3862 73922 3890
rect 78088 3884 78338 3890
rect 78036 3878 78338 3884
rect 78048 3862 78338 3878
rect 83568 3874 83858 3890
rect 94608 3874 94898 3890
rect 133248 3874 133538 3890
rect 83556 3868 83858 3874
rect 73618 3839 73674 3848
rect 59728 3810 59780 3816
rect 83608 3862 83858 3868
rect 94596 3868 94898 3874
rect 83556 3810 83608 3816
rect 94648 3862 94898 3868
rect 122288 3868 122340 3874
rect 94596 3810 94648 3816
rect 122288 3810 122340 3816
rect 133236 3868 133538 3874
rect 133288 3862 133538 3868
rect 133236 3810 133288 3816
rect 58808 3732 58860 3738
rect 58808 3674 58860 3680
rect 56048 3528 56100 3534
rect 56048 3470 56100 3476
rect 54944 3460 54996 3466
rect 54944 3402 54996 3408
rect 51356 3392 51408 3398
rect 51356 3334 51408 3340
rect 50160 3256 50212 3262
rect 50160 3198 50212 3204
rect 40960 3188 41012 3194
rect 40960 3130 41012 3136
rect 4068 1080 4120 1086
rect 4068 1022 4120 1028
rect 1676 944 1728 950
rect 1676 886 1728 892
rect 1688 480 1716 886
rect 4080 480 4108 1022
rect 19432 876 19484 882
rect 19432 818 19484 824
rect 18236 808 18288 814
rect 18236 750 18288 756
rect 9956 740 10008 746
rect 9956 682 10008 688
rect 8760 672 8812 678
rect 8760 614 8812 620
rect 8772 480 8800 614
rect 9968 480 9996 682
rect 14740 604 14792 610
rect 14740 546 14792 552
rect 17040 604 17092 610
rect 17040 546 17092 552
rect 12162 504 12218 513
rect 542 82 654 480
rect 400 66 654 82
rect 388 60 654 66
rect 440 54 654 60
rect 388 2 440 8
rect 542 -960 654 54
rect 1646 -960 1758 480
rect 2842 354 2954 480
rect 2842 338 3280 354
rect 2842 332 3292 338
rect 2842 326 3240 332
rect 2842 -960 2954 326
rect 3240 274 3292 280
rect 4038 -960 4150 480
rect 5234 354 5346 480
rect 5446 368 5502 377
rect 5234 326 5446 354
rect 5234 -960 5346 326
rect 5446 303 5502 312
rect 6274 96 6330 105
rect 6430 82 6542 480
rect 6330 54 6542 82
rect 6274 31 6330 40
rect 6430 -960 6542 54
rect 7626 218 7738 480
rect 7626 202 8064 218
rect 7626 196 8076 202
rect 7626 190 8024 196
rect 7626 -960 7738 190
rect 8024 138 8076 144
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 354 11234 480
rect 14752 480 14780 546
rect 17052 480 17080 546
rect 18248 480 18276 750
rect 19444 480 19472 818
rect 12162 439 12218 448
rect 11520 400 11572 406
rect 11122 348 11520 354
rect 11122 342 11572 348
rect 12176 354 12204 439
rect 12318 354 12430 480
rect 11122 326 11560 342
rect 12176 326 12430 354
rect 11122 -960 11234 326
rect 12318 -960 12430 326
rect 13514 218 13626 480
rect 13726 232 13782 241
rect 13514 190 13726 218
rect 13514 -960 13626 190
rect 13726 167 13782 176
rect 14710 -960 14822 480
rect 15906 354 16018 480
rect 16212 468 16264 474
rect 16212 410 16264 416
rect 16224 354 16252 410
rect 15906 326 16252 354
rect 15906 -960 16018 326
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 19812 66 19840 3060
rect 20628 1012 20680 1018
rect 20628 954 20680 960
rect 20640 480 20668 954
rect 20916 950 20944 3060
rect 20904 944 20956 950
rect 20904 886 20956 892
rect 19800 60 19852 66
rect 19800 2 19852 8
rect 20598 -960 20710 480
rect 21794 82 21906 480
rect 22020 338 22048 3060
rect 23124 1086 23152 3060
rect 23952 3046 24242 3074
rect 25056 3046 25346 3074
rect 26344 3046 26450 3074
rect 23112 1080 23164 1086
rect 23112 1022 23164 1028
rect 22008 332 22060 338
rect 22008 274 22060 280
rect 22836 264 22888 270
rect 22990 218 23102 480
rect 23952 377 23980 3046
rect 23938 368 23994 377
rect 23938 303 23994 312
rect 22888 212 23102 218
rect 22836 206 23102 212
rect 22848 190 23102 206
rect 22008 128 22060 134
rect 21794 76 22008 82
rect 21794 70 22060 76
rect 21794 54 22048 70
rect 21794 -960 21906 54
rect 22990 -960 23102 190
rect 24186 82 24298 480
rect 25056 105 25084 3046
rect 25290 354 25402 480
rect 25686 368 25742 377
rect 25290 326 25686 354
rect 25042 96 25098 105
rect 24186 66 24624 82
rect 24186 60 24636 66
rect 24186 54 24584 60
rect 24186 -960 24298 54
rect 25042 31 25098 40
rect 24584 2 24636 8
rect 25290 -960 25402 326
rect 25686 303 25742 312
rect 26344 202 26372 3046
rect 26608 2916 26660 2922
rect 26608 2858 26660 2864
rect 26620 1442 26648 2858
rect 26528 1414 26648 1442
rect 26528 480 26556 1414
rect 27540 678 27568 3060
rect 27712 2848 27764 2854
rect 27712 2790 27764 2796
rect 27528 672 27580 678
rect 27528 614 27580 620
rect 27724 480 27752 2790
rect 28644 746 28672 3060
rect 28632 740 28684 746
rect 28632 682 28684 688
rect 28906 640 28962 649
rect 28906 575 28962 584
rect 28920 480 28948 575
rect 26332 196 26384 202
rect 26332 138 26384 144
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 29748 406 29776 3060
rect 30852 513 30880 3060
rect 30838 504 30894 513
rect 29736 400 29788 406
rect 29736 342 29788 348
rect 30074 354 30186 480
rect 30838 439 30894 448
rect 30074 338 30328 354
rect 30074 332 30340 338
rect 30074 326 30288 332
rect 30074 -960 30186 326
rect 30288 274 30340 280
rect 31270 218 31382 480
rect 31956 241 31984 3060
rect 33060 542 33088 3060
rect 33600 2984 33652 2990
rect 33600 2926 33652 2932
rect 33048 536 33100 542
rect 32220 400 32272 406
rect 32374 354 32486 480
rect 33048 478 33100 484
rect 33612 480 33640 2926
rect 32272 348 32486 354
rect 32220 342 32486 348
rect 32232 326 32486 342
rect 31128 202 31382 218
rect 31116 196 31382 202
rect 31168 190 31382 196
rect 31116 138 31168 144
rect 31270 -960 31382 190
rect 31942 232 31998 241
rect 31942 167 31998 176
rect 32374 -960 32486 326
rect 33570 -960 33682 480
rect 34164 474 34192 3060
rect 34796 672 34848 678
rect 34796 614 34848 620
rect 34808 480 34836 614
rect 35268 610 35296 3060
rect 36372 814 36400 3060
rect 37476 882 37504 3060
rect 38580 1018 38608 3060
rect 39408 3046 39698 3074
rect 40512 3046 40802 3074
rect 38568 1012 38620 1018
rect 38568 954 38620 960
rect 37464 876 37516 882
rect 37464 818 37516 824
rect 36360 808 36412 814
rect 36360 750 36412 756
rect 35256 604 35308 610
rect 35256 546 35308 552
rect 35992 604 36044 610
rect 35992 546 36044 552
rect 36004 480 36032 546
rect 34152 468 34204 474
rect 34152 410 34204 416
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37002 232 37058 241
rect 37158 218 37270 480
rect 37058 190 37270 218
rect 37002 167 37058 176
rect 37158 -960 37270 190
rect 38354 354 38466 480
rect 38568 468 38620 474
rect 38568 410 38620 416
rect 38580 354 38608 410
rect 38354 326 38608 354
rect 38354 -960 38466 326
rect 39408 134 39436 3046
rect 39592 598 39804 626
rect 39592 480 39620 598
rect 39776 542 39804 598
rect 39764 536 39816 542
rect 39396 128 39448 134
rect 39396 70 39448 76
rect 39550 -960 39662 480
rect 39764 478 39816 484
rect 40512 270 40540 3046
rect 40972 1578 41000 3130
rect 40696 1550 41000 1578
rect 41616 3046 41906 3074
rect 42812 3046 43010 3074
rect 43824 3046 44114 3074
rect 44272 3052 44324 3058
rect 40696 480 40724 1550
rect 40500 264 40552 270
rect 40500 206 40552 212
rect 40654 -960 40766 480
rect 41616 66 41644 3046
rect 41850 218 41962 480
rect 42706 368 42762 377
rect 42812 354 42840 3046
rect 43824 2922 43852 3046
rect 44272 2994 44324 3000
rect 43812 2916 43864 2922
rect 43812 2858 43864 2864
rect 44284 480 44312 2994
rect 45204 2854 45232 3060
rect 45192 2848 45244 2854
rect 45192 2790 45244 2796
rect 46308 649 46336 3060
rect 46294 640 46350 649
rect 46294 575 46350 584
rect 42762 326 42840 354
rect 42706 303 42762 312
rect 42248 264 42300 270
rect 41850 212 42248 218
rect 41850 206 42300 212
rect 41850 190 42288 206
rect 41604 60 41656 66
rect 41604 2 41656 8
rect 41850 -960 41962 190
rect 43046 82 43158 480
rect 42904 66 43158 82
rect 42892 60 43158 66
rect 42944 54 43158 60
rect 42892 2 42944 8
rect 43046 -960 43158 54
rect 44242 -960 44354 480
rect 45284 128 45336 134
rect 45438 82 45550 480
rect 45336 76 45550 82
rect 45284 70 45550 76
rect 45296 54 45550 70
rect 45438 -960 45550 54
rect 46634 82 46746 480
rect 47412 338 47440 3060
rect 47860 2848 47912 2854
rect 47860 2790 47912 2796
rect 47872 480 47900 2790
rect 47400 332 47452 338
rect 47400 274 47452 280
rect 46846 96 46902 105
rect 46634 54 46846 82
rect 46634 -960 46746 54
rect 46846 31 46902 40
rect 47830 -960 47942 480
rect 48516 202 48544 3060
rect 48964 2916 49016 2922
rect 48964 2858 49016 2864
rect 48976 480 49004 2858
rect 48504 196 48556 202
rect 48504 138 48556 144
rect 48934 -960 49046 480
rect 49620 406 49648 3060
rect 50172 480 50200 3198
rect 50448 3046 50738 3074
rect 50448 2990 50476 3046
rect 50436 2984 50488 2990
rect 50436 2926 50488 2932
rect 51368 480 51396 3334
rect 52552 3120 52604 3126
rect 52552 3062 52604 3068
rect 51828 678 51856 3060
rect 51816 672 51868 678
rect 51816 614 51868 620
rect 52564 480 52592 3062
rect 52932 610 52960 3060
rect 52920 604 52972 610
rect 52920 546 52972 552
rect 49608 400 49660 406
rect 49608 342 49660 348
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 218 53830 480
rect 54036 241 54064 3060
rect 54956 480 54984 3402
rect 53576 202 53830 218
rect 53564 196 53830 202
rect 53616 190 53830 196
rect 53564 138 53616 144
rect 53718 -960 53830 190
rect 54022 232 54078 241
rect 54022 167 54078 176
rect 54914 -960 55026 480
rect 55140 474 55168 3060
rect 56060 480 56088 3470
rect 57072 3194 57362 3210
rect 57060 3188 57362 3194
rect 57112 3182 57362 3188
rect 57520 3188 57572 3194
rect 57060 3130 57112 3136
rect 57520 3130 57572 3136
rect 56244 542 56272 3060
rect 57532 1578 57560 3130
rect 57256 1550 57560 1578
rect 58176 3046 58466 3074
rect 56232 536 56284 542
rect 55128 468 55180 474
rect 55128 410 55180 416
rect 56018 -960 56130 480
rect 56232 478 56284 484
rect 57256 480 57284 1550
rect 57214 -960 57326 480
rect 58176 270 58204 3046
rect 58410 354 58522 480
rect 58820 354 58848 3674
rect 58410 326 58848 354
rect 59372 3046 59570 3074
rect 58164 264 58216 270
rect 58164 206 58216 212
rect 58410 -960 58522 326
rect 59372 66 59400 3046
rect 59740 1986 59768 3810
rect 62028 3800 62080 3806
rect 62028 3742 62080 3748
rect 67456 3800 67508 3806
rect 80888 3800 80940 3806
rect 67456 3742 67508 3748
rect 60384 3058 60674 3074
rect 60372 3052 60674 3058
rect 60424 3046 60674 3052
rect 60372 2994 60424 3000
rect 60832 2848 60884 2854
rect 60832 2790 60884 2796
rect 59648 1958 59768 1986
rect 59648 480 59676 1958
rect 60844 480 60872 2790
rect 59360 60 59412 66
rect 59360 2 59412 8
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61764 134 61792 3060
rect 62040 480 62068 3742
rect 63224 3664 63276 3670
rect 63224 3606 63276 3612
rect 61752 128 61804 134
rect 61752 70 61804 76
rect 61998 -960 62110 480
rect 62868 105 62896 3060
rect 63236 480 63264 3606
rect 66720 3596 66772 3602
rect 66720 3538 66772 3544
rect 65524 3324 65576 3330
rect 65524 3266 65576 3272
rect 63696 3046 63986 3074
rect 64328 3052 64380 3058
rect 63696 2922 63724 3046
rect 64328 2994 64380 3000
rect 64892 3046 65090 3074
rect 63684 2916 63736 2922
rect 63684 2858 63736 2864
rect 64340 480 64368 2994
rect 64892 2990 64920 3046
rect 64880 2984 64932 2990
rect 64880 2926 64932 2932
rect 65536 480 65564 3266
rect 65892 3256 65944 3262
rect 65944 3204 66194 3210
rect 65892 3198 66194 3204
rect 65904 3182 66194 3198
rect 66732 480 66760 3538
rect 67468 3398 67496 3742
rect 71424 3738 71714 3754
rect 84476 3800 84528 3806
rect 80888 3742 80940 3748
rect 69020 3732 69072 3738
rect 69020 3674 69072 3680
rect 71412 3732 71714 3738
rect 71464 3726 71714 3732
rect 71412 3674 71464 3680
rect 69032 3534 69060 3674
rect 69112 3664 69164 3670
rect 69112 3606 69164 3612
rect 69020 3528 69072 3534
rect 69020 3470 69072 3476
rect 66996 3392 67048 3398
rect 67456 3392 67508 3398
rect 67048 3340 67298 3346
rect 66996 3334 67298 3340
rect 67456 3334 67508 3340
rect 67008 3318 67298 3334
rect 68100 3120 68152 3126
rect 68152 3068 68402 3074
rect 68100 3062 68402 3068
rect 68112 3046 68402 3062
rect 67916 2984 67968 2990
rect 67916 2926 67968 2932
rect 67928 480 67956 2926
rect 69124 480 69152 3606
rect 70124 3528 70176 3534
rect 70124 3470 70176 3476
rect 72976 3528 73028 3534
rect 72976 3470 73028 3476
rect 78588 3528 78640 3534
rect 78588 3470 78640 3476
rect 62854 96 62910 105
rect 62854 31 62910 40
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 69492 202 69520 3060
rect 70136 218 70164 3470
rect 70216 3460 70268 3466
rect 70216 3402 70268 3408
rect 70228 3346 70256 3402
rect 70228 3318 70610 3346
rect 71504 3324 71556 3330
rect 71504 3266 71556 3272
rect 71516 480 71544 3266
rect 72528 3194 72818 3210
rect 72516 3188 72818 3194
rect 72568 3182 72818 3188
rect 72516 3130 72568 3136
rect 70278 218 70390 480
rect 69480 196 69532 202
rect 70136 190 70390 218
rect 69480 138 69532 144
rect 70278 -960 70390 190
rect 71474 -960 71586 480
rect 72578 354 72690 480
rect 72988 354 73016 3470
rect 76932 3392 76984 3398
rect 76984 3340 77234 3346
rect 76932 3334 77234 3340
rect 76944 3318 77234 3334
rect 73804 3188 73856 3194
rect 73804 3130 73856 3136
rect 73816 480 73844 3130
rect 76288 3120 76340 3126
rect 75840 3046 76130 3074
rect 76288 3062 76340 3068
rect 75368 2916 75420 2922
rect 75368 2858 75420 2864
rect 72578 326 73016 354
rect 72578 -960 72690 326
rect 73774 -960 73886 480
rect 74970 354 75082 480
rect 75380 354 75408 2858
rect 75840 2854 75868 3046
rect 75828 2848 75880 2854
rect 75828 2790 75880 2796
rect 76300 1578 76328 3062
rect 77392 2848 77444 2854
rect 77392 2790 77444 2796
rect 76208 1550 76328 1578
rect 76208 480 76236 1550
rect 77404 480 77432 2790
rect 78600 480 78628 3470
rect 79692 3392 79744 3398
rect 79692 3334 79744 3340
rect 79600 3120 79652 3126
rect 79152 3058 79442 3074
rect 79600 3062 79652 3068
rect 79140 3052 79442 3058
rect 79192 3046 79442 3052
rect 79140 2994 79192 3000
rect 79612 2922 79640 3062
rect 79600 2916 79652 2922
rect 79600 2858 79652 2864
rect 79704 480 79732 3334
rect 79968 3256 80020 3262
rect 80020 3204 80546 3210
rect 79968 3198 80546 3204
rect 79980 3182 80546 3198
rect 80900 480 80928 3742
rect 81360 3738 81650 3754
rect 84476 3742 84528 3748
rect 98000 3800 98052 3806
rect 114008 3800 114060 3806
rect 98052 3748 98210 3754
rect 98000 3742 98210 3748
rect 81348 3732 81650 3738
rect 81400 3726 81650 3732
rect 81348 3674 81400 3680
rect 82912 3596 82964 3602
rect 82912 3538 82964 3544
rect 83280 3596 83332 3602
rect 83280 3538 83332 3544
rect 82924 3330 82952 3538
rect 83004 3392 83056 3398
rect 83004 3334 83056 3340
rect 82912 3324 82964 3330
rect 82912 3266 82964 3272
rect 82740 2990 82768 3060
rect 83016 3058 83044 3334
rect 83004 3052 83056 3058
rect 83004 2994 83056 3000
rect 82728 2984 82780 2990
rect 82728 2926 82780 2932
rect 82084 2916 82136 2922
rect 82084 2858 82136 2864
rect 82096 480 82124 2858
rect 83292 480 83320 3538
rect 84488 480 84516 3742
rect 85672 3732 85724 3738
rect 85672 3674 85724 3680
rect 87788 3732 87840 3738
rect 98012 3726 98210 3742
rect 101232 3738 101522 3754
rect 114008 3742 114060 3748
rect 101220 3732 101522 3738
rect 87788 3674 87840 3680
rect 101272 3726 101522 3732
rect 101220 3674 101272 3680
rect 84672 3330 84962 3346
rect 84660 3324 84962 3330
rect 84712 3318 84962 3324
rect 84660 3266 84712 3272
rect 85684 480 85712 3674
rect 86868 3664 86920 3670
rect 86920 3612 87170 3618
rect 86868 3606 87170 3612
rect 86880 3590 87170 3606
rect 85776 3466 86066 3482
rect 85764 3460 86066 3466
rect 85816 3454 86066 3460
rect 85764 3402 85816 3408
rect 86868 3324 86920 3330
rect 86868 3266 86920 3272
rect 86880 480 86908 3266
rect 74970 326 75408 354
rect 74970 -960 75082 326
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87800 218 87828 3674
rect 99012 3664 99064 3670
rect 96816 3602 97106 3618
rect 109408 3664 109460 3670
rect 99064 3612 99314 3618
rect 99012 3606 99314 3612
rect 109408 3606 109460 3612
rect 96804 3596 97106 3602
rect 96856 3590 97106 3596
rect 99024 3590 99314 3606
rect 102232 3596 102284 3602
rect 96804 3538 96856 3544
rect 102232 3538 102284 3544
rect 92388 3528 92440 3534
rect 92440 3476 92690 3482
rect 92388 3470 92690 3476
rect 90364 3460 90416 3466
rect 92400 3454 92690 3470
rect 90364 3402 90416 3408
rect 89536 3392 89588 3398
rect 89536 3334 89588 3340
rect 87984 3194 88274 3210
rect 87972 3188 88274 3194
rect 88024 3182 88274 3188
rect 87972 3130 88024 3136
rect 89076 3120 89128 3126
rect 89128 3068 89378 3074
rect 89076 3062 89378 3068
rect 89088 3046 89378 3062
rect 87942 218 88054 480
rect 87800 190 88054 218
rect 87942 -960 88054 190
rect 89138 354 89250 480
rect 89548 354 89576 3334
rect 90376 480 90404 3402
rect 96252 3392 96304 3398
rect 96252 3334 96304 3340
rect 93952 3256 94004 3262
rect 93952 3198 94004 3204
rect 90468 2990 90496 3060
rect 91296 3046 91586 3074
rect 93504 3058 93794 3074
rect 93492 3052 93794 3058
rect 90456 2984 90508 2990
rect 90456 2926 90508 2932
rect 91296 2854 91324 3046
rect 93544 3046 93794 3052
rect 93492 2994 93544 3000
rect 91560 2984 91612 2990
rect 91560 2926 91612 2932
rect 91284 2848 91336 2854
rect 91284 2790 91336 2796
rect 91572 480 91600 2926
rect 92756 2848 92808 2854
rect 92756 2790 92808 2796
rect 92768 480 92796 2790
rect 93964 480 93992 3198
rect 95148 3052 95200 3058
rect 95148 2994 95200 3000
rect 95160 480 95188 2994
rect 95988 2922 96016 3060
rect 95976 2916 96028 2922
rect 95976 2858 96028 2864
rect 96264 480 96292 3334
rect 100128 3330 100418 3346
rect 100116 3324 100418 3330
rect 100168 3318 100418 3324
rect 100116 3266 100168 3272
rect 101036 3188 101088 3194
rect 101036 3130 101088 3136
rect 98736 3120 98788 3126
rect 98736 3062 98788 3068
rect 97448 2916 97500 2922
rect 97448 2858 97500 2864
rect 97460 480 97488 2858
rect 98644 2848 98696 2854
rect 98644 2790 98696 2796
rect 98656 1290 98684 2790
rect 98644 1284 98696 1290
rect 98644 1226 98696 1232
rect 98748 1170 98776 3062
rect 99840 2848 99892 2854
rect 99840 2790 99892 2796
rect 98656 1142 98776 1170
rect 98656 480 98684 1142
rect 99852 480 99880 2790
rect 101048 480 101076 3130
rect 102244 480 102272 3538
rect 103612 3528 103664 3534
rect 102336 3466 102626 3482
rect 103664 3476 103730 3482
rect 103612 3470 103730 3476
rect 102324 3460 102626 3466
rect 102376 3454 102626 3460
rect 103624 3454 103730 3470
rect 105728 3460 105780 3466
rect 102324 3402 102376 3408
rect 105728 3402 105780 3408
rect 103336 3324 103388 3330
rect 103336 3266 103388 3272
rect 103348 480 103376 3266
rect 104544 3046 104834 3074
rect 104544 2990 104572 3046
rect 104532 2984 104584 2990
rect 104532 2926 104584 2932
rect 104624 2984 104676 2990
rect 104624 2926 104676 2932
rect 104636 1578 104664 2926
rect 104544 1550 104664 1578
rect 104544 480 104572 1550
rect 105740 480 105768 3402
rect 109040 3392 109092 3398
rect 109092 3340 109250 3346
rect 109040 3334 109250 3340
rect 109052 3318 109250 3334
rect 106740 3256 106792 3262
rect 107200 3256 107252 3262
rect 106792 3204 107042 3210
rect 106740 3198 107042 3204
rect 107200 3198 107252 3204
rect 106752 3182 107042 3198
rect 105924 1290 105952 3060
rect 107212 1714 107240 3198
rect 107856 3058 108146 3074
rect 107844 3052 108146 3058
rect 107896 3046 108146 3052
rect 108488 3052 108540 3058
rect 107844 2994 107896 3000
rect 108488 2994 108540 3000
rect 106936 1686 107240 1714
rect 105912 1284 105964 1290
rect 105912 1226 105964 1232
rect 106936 480 106964 1686
rect 89138 326 89576 354
rect 89138 -960 89250 326
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 354 108202 480
rect 108500 354 108528 2994
rect 109420 1850 109448 3606
rect 110512 3528 110564 3534
rect 110512 3470 110564 3476
rect 110064 3046 110354 3074
rect 110064 2922 110092 3046
rect 110052 2916 110104 2922
rect 110052 2858 110104 2864
rect 109328 1822 109448 1850
rect 109328 480 109356 1822
rect 110524 480 110552 3470
rect 112812 3392 112864 3398
rect 112812 3334 112864 3340
rect 111156 3120 111208 3126
rect 111616 3120 111668 3126
rect 111208 3068 111458 3074
rect 111156 3062 111458 3068
rect 111616 3062 111668 3068
rect 111168 3046 111458 3062
rect 111628 480 111656 3062
rect 112548 2854 112576 3060
rect 112536 2848 112588 2854
rect 112536 2790 112588 2796
rect 112824 480 112852 3334
rect 113100 3194 113666 3210
rect 113088 3188 113666 3194
rect 113140 3182 113666 3188
rect 113088 3130 113140 3136
rect 114020 480 114048 3742
rect 116400 3732 116452 3738
rect 116400 3674 116452 3680
rect 114480 3602 114770 3618
rect 114468 3596 114770 3602
rect 114520 3590 114770 3596
rect 114468 3538 114520 3544
rect 115584 3330 115874 3346
rect 115572 3324 115874 3330
rect 115624 3318 115874 3324
rect 115572 3266 115624 3272
rect 115204 2916 115256 2922
rect 115204 2858 115256 2864
rect 115216 480 115244 2858
rect 116412 480 116440 3674
rect 121184 3664 121236 3670
rect 121236 3612 121394 3618
rect 121184 3606 121394 3612
rect 121092 3596 121144 3602
rect 121196 3590 121394 3606
rect 121092 3538 121144 3544
rect 117792 3466 118082 3482
rect 117780 3460 118082 3466
rect 117832 3454 118082 3460
rect 117780 3402 117832 3408
rect 117596 3324 117648 3330
rect 117596 3266 117648 3272
rect 116964 2990 116992 3060
rect 116952 2984 117004 2990
rect 116952 2926 117004 2932
rect 117608 480 117636 3266
rect 118608 3256 118660 3262
rect 119896 3256 119948 3262
rect 118660 3204 119186 3210
rect 118608 3198 119186 3204
rect 119896 3198 119948 3204
rect 118620 3182 119186 3198
rect 118792 2848 118844 2854
rect 118792 2790 118844 2796
rect 118804 480 118832 2790
rect 119908 480 119936 3198
rect 120000 3058 120290 3074
rect 119988 3052 120290 3058
rect 120040 3046 120290 3052
rect 119988 2994 120040 3000
rect 121104 480 121132 3538
rect 122300 480 122328 3810
rect 125508 3800 125560 3806
rect 125560 3748 125810 3754
rect 125508 3742 125810 3748
rect 125520 3726 125810 3742
rect 127728 3738 128018 3754
rect 127716 3732 128018 3738
rect 127768 3726 128018 3732
rect 127716 3674 127768 3680
rect 125048 3664 125100 3670
rect 135444 3664 135496 3670
rect 125048 3606 125100 3612
rect 122380 3528 122432 3534
rect 122432 3476 122498 3482
rect 122380 3470 122498 3476
rect 122392 3454 122498 3470
rect 124128 3392 124180 3398
rect 124180 3340 124706 3346
rect 124128 3334 124706 3340
rect 124140 3318 124706 3334
rect 123300 3120 123352 3126
rect 123352 3068 123602 3074
rect 123300 3062 123602 3068
rect 123312 3046 123602 3062
rect 123484 2984 123536 2990
rect 123484 2926 123536 2932
rect 123496 480 123524 2926
rect 108090 326 108528 354
rect 108090 -960 108202 326
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 354 124762 480
rect 125060 354 125088 3606
rect 132144 3602 132434 3618
rect 143632 3664 143684 3670
rect 135496 3612 135746 3618
rect 135444 3606 135746 3612
rect 153108 3664 153160 3670
rect 143632 3606 143684 3612
rect 132132 3596 132434 3602
rect 132184 3590 132434 3596
rect 135456 3590 135746 3606
rect 136456 3596 136508 3602
rect 132132 3538 132184 3544
rect 136456 3538 136508 3544
rect 127072 3528 127124 3534
rect 127072 3470 127124 3476
rect 125968 3392 126020 3398
rect 125968 3334 126020 3340
rect 125980 1714 126008 3334
rect 126900 2922 126928 3060
rect 126888 2916 126940 2922
rect 126888 2858 126940 2864
rect 127084 1850 127112 3470
rect 131764 3460 131816 3466
rect 131764 3402 131816 3408
rect 128832 3330 129122 3346
rect 128820 3324 129122 3330
rect 128872 3318 129122 3324
rect 129372 3324 129424 3330
rect 128820 3266 128872 3272
rect 129372 3266 129424 3272
rect 128176 3052 128228 3058
rect 128176 2994 128228 3000
rect 125888 1686 126008 1714
rect 126992 1822 127112 1850
rect 125888 480 125916 1686
rect 126992 480 127020 1822
rect 128188 480 128216 2994
rect 129384 480 129412 3266
rect 131028 3256 131080 3262
rect 131080 3204 131330 3210
rect 131028 3198 131330 3204
rect 131040 3182 131330 3198
rect 130212 2854 130240 3060
rect 130568 2984 130620 2990
rect 130568 2926 130620 2932
rect 130200 2848 130252 2854
rect 130200 2790 130252 2796
rect 130580 480 130608 2926
rect 131776 480 131804 3402
rect 134352 3194 134642 3210
rect 134340 3188 134642 3194
rect 134392 3182 134642 3188
rect 134340 3130 134392 3136
rect 134156 3120 134208 3126
rect 134156 3062 134208 3068
rect 132960 2916 133012 2922
rect 132960 2858 133012 2864
rect 132972 480 133000 2858
rect 134168 480 134196 3062
rect 135260 2848 135312 2854
rect 135260 2790 135312 2796
rect 135272 480 135300 2790
rect 136468 480 136496 3538
rect 137652 3528 137704 3534
rect 139216 3528 139268 3534
rect 137704 3476 137954 3482
rect 137652 3470 137954 3476
rect 139216 3470 139268 3476
rect 137664 3454 137954 3470
rect 136640 3392 136692 3398
rect 136692 3340 136850 3346
rect 136640 3334 136850 3340
rect 136652 3318 136850 3334
rect 137652 3188 137704 3194
rect 137652 3130 137704 3136
rect 137664 480 137692 3130
rect 138768 3058 139058 3074
rect 138756 3052 139058 3058
rect 138808 3046 139058 3052
rect 138756 2994 138808 3000
rect 124650 326 125088 354
rect 124650 -960 124762 326
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 354 138930 480
rect 139228 354 139256 3470
rect 142264 3466 142370 3482
rect 142252 3460 142370 3466
rect 142304 3454 142370 3460
rect 142528 3460 142580 3466
rect 142252 3402 142304 3408
rect 142528 3402 142580 3408
rect 139872 3330 140162 3346
rect 139860 3324 140162 3330
rect 139912 3318 140162 3324
rect 139860 3266 139912 3272
rect 140044 3256 140096 3262
rect 140044 3198 140096 3204
rect 140056 480 140084 3198
rect 140976 3046 141266 3074
rect 140976 2990 141004 3046
rect 140964 2984 141016 2990
rect 140964 2926 141016 2932
rect 141240 2984 141292 2990
rect 141240 2926 141292 2932
rect 141252 480 141280 2926
rect 142540 1578 142568 3402
rect 143184 3058 143474 3074
rect 143172 3052 143474 3058
rect 143224 3046 143474 3052
rect 143172 2994 143224 3000
rect 143644 1850 143672 3606
rect 146496 3602 146786 3618
rect 153160 3612 153410 3618
rect 153108 3606 153410 3612
rect 146484 3596 146786 3602
rect 146536 3590 146786 3596
rect 149520 3596 149572 3602
rect 146484 3538 146536 3544
rect 153120 3590 153410 3606
rect 158640 3602 158930 3618
rect 158628 3596 158930 3602
rect 149520 3538 149572 3544
rect 158680 3590 158930 3596
rect 158628 3538 158680 3544
rect 148692 3528 148744 3534
rect 148744 3476 148994 3482
rect 148692 3470 148994 3476
rect 148704 3454 148994 3470
rect 148324 3324 148376 3330
rect 148324 3266 148376 3272
rect 147784 3194 147890 3210
rect 147772 3188 147890 3194
rect 147824 3182 147890 3188
rect 147772 3130 147824 3136
rect 144276 3120 144328 3126
rect 147128 3120 147180 3126
rect 144328 3068 144578 3074
rect 144276 3062 144578 3068
rect 144288 3046 144578 3062
rect 145392 3046 145682 3074
rect 147128 3062 147180 3068
rect 145932 3052 145984 3058
rect 144736 2916 144788 2922
rect 144736 2858 144788 2864
rect 142448 1550 142568 1578
rect 143552 1822 143672 1850
rect 142448 480 142476 1550
rect 143552 480 143580 1822
rect 144748 480 144776 2858
rect 145392 2854 145420 3046
rect 145932 2994 145984 3000
rect 145380 2848 145432 2854
rect 145380 2790 145432 2796
rect 145944 480 145972 2994
rect 147140 480 147168 3062
rect 148336 480 148364 3266
rect 149532 480 149560 3538
rect 153016 3528 153068 3534
rect 151740 3466 152306 3482
rect 153016 3470 153068 3476
rect 160192 3528 160244 3534
rect 160192 3470 160244 3476
rect 151728 3460 152306 3466
rect 151780 3454 152306 3460
rect 151728 3402 151780 3408
rect 149796 3392 149848 3398
rect 149848 3340 150098 3346
rect 149796 3334 150098 3340
rect 149808 3318 150098 3334
rect 150912 3046 151202 3074
rect 151820 3052 151872 3058
rect 150912 2990 150940 3046
rect 151820 2994 151872 3000
rect 150900 2984 150952 2990
rect 150900 2926 150952 2932
rect 150624 2916 150676 2922
rect 150624 2858 150676 2864
rect 150636 480 150664 2858
rect 151832 480 151860 2994
rect 153028 480 153056 3470
rect 155776 3460 155828 3466
rect 155776 3402 155828 3408
rect 154028 3256 154080 3262
rect 154028 3198 154080 3204
rect 138818 326 139256 354
rect 138818 -960 138930 326
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154040 218 154068 3198
rect 155316 3120 155368 3126
rect 154224 3046 154514 3074
rect 155368 3068 155618 3074
rect 155316 3062 155618 3068
rect 155328 3046 155618 3062
rect 154224 2854 154252 3046
rect 154212 2848 154264 2854
rect 154212 2790 154264 2796
rect 154182 218 154294 480
rect 154040 190 154294 218
rect 154182 -960 154294 190
rect 155378 354 155490 480
rect 155788 354 155816 3402
rect 157260 3330 157826 3346
rect 157248 3324 157826 3330
rect 157300 3318 157826 3324
rect 158168 3324 158220 3330
rect 157248 3266 157300 3272
rect 158168 3266 158220 3272
rect 156432 3194 156722 3210
rect 156420 3188 156722 3194
rect 156472 3182 156722 3188
rect 156420 3130 156472 3136
rect 156604 2984 156656 2990
rect 156604 2926 156656 2932
rect 156616 480 156644 2926
rect 155378 326 155816 354
rect 155378 -960 155490 326
rect 156574 -960 156686 480
rect 157770 354 157882 480
rect 158180 354 158208 3266
rect 160204 3262 160232 3470
rect 166080 3460 166132 3466
rect 166080 3402 166132 3408
rect 161296 3324 161348 3330
rect 161296 3266 161348 3272
rect 160192 3256 160244 3262
rect 160192 3198 160244 3204
rect 160020 2922 160048 3060
rect 160848 3058 161138 3074
rect 160836 3052 161138 3058
rect 160888 3046 161138 3052
rect 160836 2994 160888 3000
rect 160008 2916 160060 2922
rect 160008 2858 160060 2864
rect 160100 2916 160152 2922
rect 160100 2858 160152 2864
rect 158904 2848 158956 2854
rect 158904 2790 158956 2796
rect 158916 480 158944 2790
rect 160112 480 160140 2858
rect 161308 480 161336 3266
rect 161940 3256 161992 3262
rect 163688 3256 163740 3262
rect 161992 3204 162242 3210
rect 161940 3198 162242 3204
rect 163688 3198 163740 3204
rect 161952 3182 162242 3198
rect 162768 3120 162820 3126
rect 162820 3068 163346 3074
rect 162768 3062 163346 3068
rect 162492 3052 162544 3058
rect 162780 3046 163346 3062
rect 162492 2994 162544 3000
rect 162504 480 162532 2994
rect 163700 480 163728 3198
rect 164160 3194 164450 3210
rect 164148 3188 164450 3194
rect 164200 3182 164450 3188
rect 164148 3130 164200 3136
rect 164884 3120 164936 3126
rect 164884 3062 164936 3068
rect 164896 480 164924 3062
rect 165540 2990 165568 3060
rect 165528 2984 165580 2990
rect 165528 2926 165580 2932
rect 166092 480 166120 3402
rect 166356 3392 166408 3398
rect 174084 3392 174136 3398
rect 166408 3340 166658 3346
rect 166356 3334 166658 3340
rect 166368 3318 166658 3334
rect 169680 3330 169970 3346
rect 174136 3340 174386 3346
rect 174084 3334 174386 3340
rect 169668 3324 169970 3330
rect 169720 3318 169970 3324
rect 174096 3318 174386 3334
rect 181824 3330 182114 3346
rect 181812 3324 182114 3330
rect 169668 3266 169720 3272
rect 181864 3318 182114 3324
rect 564190 3330 564388 3346
rect 564190 3324 564400 3330
rect 564190 3318 564348 3324
rect 181812 3266 181864 3272
rect 564348 3266 564400 3272
rect 583392 3324 583444 3330
rect 583392 3266 583444 3272
rect 171876 3256 171928 3262
rect 174268 3256 174320 3262
rect 171928 3204 172178 3210
rect 171876 3198 172178 3204
rect 180892 3256 180944 3262
rect 174268 3198 174320 3204
rect 170772 3188 170824 3194
rect 171888 3182 172178 3198
rect 170772 3130 170824 3136
rect 167184 2984 167236 2990
rect 167184 2926 167236 2932
rect 167196 480 167224 2926
rect 167748 2854 167776 3060
rect 168852 2922 168880 3060
rect 168840 2916 168892 2922
rect 168840 2858 168892 2864
rect 169576 2916 169628 2922
rect 169576 2858 169628 2864
rect 167736 2848 167788 2854
rect 167736 2790 167788 2796
rect 168380 2848 168432 2854
rect 168380 2790 168432 2796
rect 168392 480 168420 2790
rect 169588 480 169616 2858
rect 170784 480 170812 3130
rect 172980 3120 173032 3126
rect 170876 3058 171074 3074
rect 173440 3120 173492 3126
rect 173032 3068 173282 3074
rect 172980 3062 173282 3068
rect 173440 3062 173492 3068
rect 170864 3052 171074 3058
rect 170916 3046 171074 3052
rect 171968 3052 172020 3058
rect 170864 2994 170916 3000
rect 172992 3046 173282 3062
rect 171968 2994 172020 3000
rect 171980 480 172008 2994
rect 173452 1714 173480 3062
rect 173176 1686 173480 1714
rect 173176 480 173204 1686
rect 174280 480 174308 3198
rect 178512 3194 178802 3210
rect 184940 3256 184992 3262
rect 180944 3204 181010 3210
rect 180892 3198 181010 3204
rect 200304 3256 200356 3262
rect 184940 3198 184992 3204
rect 178500 3188 178802 3194
rect 178552 3182 178802 3188
rect 180904 3182 181010 3198
rect 181444 3188 181496 3194
rect 178500 3130 178552 3136
rect 181444 3130 181496 3136
rect 179052 3120 179104 3126
rect 175476 2990 175504 3060
rect 176304 3046 176594 3074
rect 179052 3062 179104 3068
rect 175464 2984 175516 2990
rect 175464 2926 175516 2932
rect 175832 2984 175884 2990
rect 175832 2926 175884 2932
rect 157770 326 158208 354
rect 157770 -960 157882 326
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 354 175546 480
rect 175844 354 175872 2926
rect 176304 2854 176332 3046
rect 177684 2922 177712 3060
rect 177856 2984 177908 2990
rect 177856 2926 177908 2932
rect 177672 2916 177724 2922
rect 177672 2858 177724 2864
rect 176292 2848 176344 2854
rect 176292 2790 176344 2796
rect 176660 1352 176712 1358
rect 176660 1294 176712 1300
rect 176672 480 176700 1294
rect 177868 480 177896 2926
rect 179064 480 179092 3062
rect 179616 3058 179906 3074
rect 179604 3052 179906 3058
rect 179656 3046 179906 3052
rect 179604 2994 179656 3000
rect 180248 2848 180300 2854
rect 180248 2790 180300 2796
rect 180260 480 180288 2790
rect 181456 480 181484 3130
rect 182548 3052 182600 3058
rect 182548 2994 182600 3000
rect 182928 3046 183218 3074
rect 182560 480 182588 2994
rect 182928 2922 182956 3046
rect 182916 2916 182968 2922
rect 182916 2858 182968 2864
rect 183744 2916 183796 2922
rect 183744 2858 183796 2864
rect 183756 480 183784 2858
rect 184308 1358 184336 3060
rect 184296 1352 184348 1358
rect 184296 1294 184348 1300
rect 184952 480 184980 3198
rect 188448 3194 188738 3210
rect 188436 3188 188738 3194
rect 188488 3182 188738 3188
rect 189552 3182 189842 3210
rect 191760 3194 192050 3210
rect 206100 3256 206152 3262
rect 200304 3198 200356 3204
rect 191748 3188 192050 3194
rect 188436 3130 188488 3136
rect 186320 3120 186372 3126
rect 186372 3068 186530 3074
rect 186320 3062 186530 3068
rect 185412 2990 185440 3060
rect 186332 3046 186530 3062
rect 187344 3046 187634 3074
rect 189552 3058 189580 3182
rect 191800 3182 192050 3188
rect 195612 3188 195664 3194
rect 191748 3130 191800 3136
rect 195612 3130 195664 3136
rect 190552 3120 190604 3126
rect 190552 3062 190604 3068
rect 189540 3052 189592 3058
rect 185400 2984 185452 2990
rect 185400 2926 185452 2932
rect 187344 2854 187372 3046
rect 189540 2994 189592 3000
rect 189724 3052 189776 3058
rect 189724 2994 189776 3000
rect 187332 2848 187384 2854
rect 187332 2790 187384 2796
rect 187332 1352 187384 1358
rect 187332 1294 187384 1300
rect 186136 1216 186188 1222
rect 186136 1158 186188 1164
rect 186148 480 186176 1158
rect 187344 480 187372 1294
rect 188896 1284 188948 1290
rect 188896 1226 188948 1232
rect 175434 326 175872 354
rect 175434 -960 175546 326
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 354 188610 480
rect 188908 354 188936 1226
rect 189736 480 189764 2994
rect 188498 326 188936 354
rect 188498 -960 188610 326
rect 189694 -960 189806 480
rect 190564 354 190592 3062
rect 190656 3046 190946 3074
rect 190656 2922 190684 3046
rect 190644 2916 190696 2922
rect 190644 2858 190696 2864
rect 192392 2916 192444 2922
rect 192392 2858 192444 2864
rect 190798 354 190910 480
rect 190564 326 190910 354
rect 190798 -960 190910 326
rect 191994 354 192106 480
rect 192404 354 192432 2858
rect 193140 1222 193168 3060
rect 193220 2780 193272 2786
rect 193220 2722 193272 2728
rect 193128 1216 193180 1222
rect 193128 1158 193180 1164
rect 193232 480 193260 2722
rect 194244 1358 194272 3060
rect 194416 2984 194468 2990
rect 194416 2926 194468 2932
rect 194232 1352 194284 1358
rect 194232 1294 194284 1300
rect 194428 480 194456 2926
rect 195348 1290 195376 3060
rect 195336 1284 195388 1290
rect 195336 1226 195388 1232
rect 195624 480 195652 3130
rect 197268 3120 197320 3126
rect 196176 3058 196466 3074
rect 197320 3068 197570 3074
rect 197268 3062 197570 3068
rect 196164 3052 196466 3058
rect 196216 3046 196466 3052
rect 197280 3046 197570 3062
rect 198384 3046 198674 3074
rect 199488 3046 199778 3074
rect 196164 2994 196216 3000
rect 198384 2922 198412 3046
rect 199108 2984 199160 2990
rect 199108 2926 199160 2932
rect 198372 2916 198424 2922
rect 198372 2858 198424 2864
rect 198280 1352 198332 1358
rect 198280 1294 198332 1300
rect 197176 1284 197228 1290
rect 197176 1226 197228 1232
rect 191994 326 192432 354
rect 191994 -960 192106 326
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 354 196890 480
rect 197188 354 197216 1226
rect 196778 326 197216 354
rect 197882 354 197994 480
rect 198292 354 198320 1294
rect 199120 480 199148 2926
rect 199488 2854 199516 3046
rect 199476 2848 199528 2854
rect 199476 2790 199528 2796
rect 200316 480 200344 3198
rect 201696 3194 201986 3210
rect 556712 3256 556764 3262
rect 206152 3204 206402 3210
rect 206100 3198 206402 3204
rect 201684 3188 201986 3194
rect 201736 3182 201986 3188
rect 206112 3182 206402 3198
rect 224880 3194 225170 3210
rect 220268 3188 220320 3194
rect 201684 3130 201736 3136
rect 220268 3130 220320 3136
rect 224868 3188 225170 3194
rect 224920 3182 225170 3188
rect 556462 3204 556712 3210
rect 575112 3256 575164 3262
rect 556462 3198 556764 3204
rect 556462 3182 556752 3198
rect 560878 3194 561168 3210
rect 575112 3198 575164 3204
rect 560878 3188 561180 3194
rect 560878 3182 561128 3188
rect 224868 3130 224920 3136
rect 561128 3130 561180 3136
rect 202696 3120 202748 3126
rect 200592 3058 200882 3074
rect 208308 3120 208360 3126
rect 202696 3062 202748 3068
rect 200580 3052 200882 3058
rect 200632 3046 200882 3052
rect 200580 2994 200632 3000
rect 201500 2916 201552 2922
rect 201500 2858 201552 2864
rect 201512 480 201540 2858
rect 202708 480 202736 3062
rect 203076 1290 203104 3060
rect 203892 3052 203944 3058
rect 203892 2994 203944 3000
rect 203064 1284 203116 1290
rect 203064 1226 203116 1232
rect 203904 480 203932 2994
rect 204180 1358 204208 3060
rect 205008 3046 205298 3074
rect 206940 3046 207506 3074
rect 209872 3120 209924 3126
rect 208360 3068 208610 3074
rect 208308 3062 208610 3068
rect 208320 3046 208610 3062
rect 209424 3058 209714 3074
rect 214932 3120 214984 3126
rect 209872 3062 209924 3068
rect 209412 3052 209714 3058
rect 205008 2990 205036 3046
rect 206940 2990 206968 3046
rect 209464 3046 209714 3052
rect 209412 2994 209464 3000
rect 204996 2984 205048 2990
rect 204996 2926 205048 2932
rect 206928 2984 206980 2990
rect 206928 2926 206980 2932
rect 208584 2984 208636 2990
rect 208584 2926 208636 2932
rect 206192 2916 206244 2922
rect 206192 2858 206244 2864
rect 205088 2848 205140 2854
rect 205088 2790 205140 2796
rect 204168 1352 204220 1358
rect 204168 1294 204220 1300
rect 205100 480 205128 2790
rect 206204 480 206232 2858
rect 207388 1352 207440 1358
rect 207388 1294 207440 1300
rect 207400 480 207428 1294
rect 208596 480 208624 2926
rect 209884 1578 209912 3062
rect 210528 3046 210818 3074
rect 211632 3046 211922 3074
rect 212172 3052 212224 3058
rect 210528 2854 210556 3046
rect 211632 2922 211660 3046
rect 212172 2994 212224 3000
rect 211620 2916 211672 2922
rect 211620 2858 211672 2864
rect 210516 2848 210568 2854
rect 210516 2790 210568 2796
rect 210976 2848 211028 2854
rect 210976 2790 211028 2796
rect 209792 1550 209912 1578
rect 209792 480 209820 1550
rect 210988 480 211016 2790
rect 212184 480 212212 2994
rect 213012 1358 213040 3060
rect 213840 3046 214130 3074
rect 215668 3120 215720 3126
rect 214984 3068 215234 3074
rect 214932 3062 215234 3068
rect 215668 3062 215720 3068
rect 214944 3046 215234 3062
rect 213840 2990 213868 3046
rect 213828 2984 213880 2990
rect 213828 2926 213880 2932
rect 214472 2984 214524 2990
rect 214472 2926 214524 2932
rect 213368 2916 213420 2922
rect 213368 2858 213420 2864
rect 213000 1352 213052 1358
rect 213000 1294 213052 1300
rect 213380 480 213408 2858
rect 214484 480 214512 2926
rect 215680 480 215708 3062
rect 216048 3046 216338 3074
rect 217152 3058 217442 3074
rect 217140 3052 217442 3058
rect 216048 2854 216076 3046
rect 217192 3046 217442 3052
rect 217980 3046 218546 3074
rect 219256 3052 219308 3058
rect 217140 2994 217192 3000
rect 217980 2922 218008 3046
rect 219256 2994 219308 3000
rect 219360 3046 219650 3074
rect 217968 2916 218020 2922
rect 217968 2858 218020 2864
rect 218060 2916 218112 2922
rect 218060 2858 218112 2864
rect 216036 2848 216088 2854
rect 216036 2790 216088 2796
rect 216864 2848 216916 2854
rect 216864 2790 216916 2796
rect 216876 480 216904 2790
rect 218072 480 218100 2858
rect 219268 480 219296 2994
rect 219360 2990 219388 3046
rect 219348 2984 219400 2990
rect 219348 2926 219400 2932
rect 197882 326 198320 354
rect 196778 -960 196890 326
rect 197882 -960 197994 326
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220280 218 220308 3130
rect 220452 3120 220504 3126
rect 221556 3120 221608 3126
rect 220504 3068 220754 3074
rect 220452 3062 220754 3068
rect 225972 3120 226024 3126
rect 221556 3062 221608 3068
rect 220464 3046 220754 3062
rect 221568 480 221596 3062
rect 221844 2854 221872 3060
rect 222948 2922 222976 3060
rect 223500 3058 224066 3074
rect 228732 3120 228784 3126
rect 226024 3068 226274 3074
rect 225972 3062 226274 3068
rect 223488 3052 224066 3058
rect 223540 3046 224066 3052
rect 225984 3046 226274 3062
rect 223488 2994 223540 3000
rect 223948 2984 224000 2990
rect 223948 2926 224000 2932
rect 225144 2984 225196 2990
rect 225144 2926 225196 2932
rect 222936 2916 222988 2922
rect 222936 2858 222988 2864
rect 223120 2916 223172 2922
rect 223120 2858 223172 2864
rect 221832 2848 221884 2854
rect 221832 2790 221884 2796
rect 220422 218 220534 480
rect 220280 190 220534 218
rect 220422 -960 220534 190
rect 221526 -960 221638 480
rect 222722 354 222834 480
rect 223132 354 223160 2858
rect 223960 480 223988 2926
rect 225156 480 225184 2926
rect 227364 2922 227392 3060
rect 228192 3058 228482 3074
rect 228732 3062 228784 3068
rect 232596 3120 232648 3126
rect 239312 3120 239364 3126
rect 232648 3068 232898 3074
rect 232596 3062 232898 3068
rect 228180 3052 228482 3058
rect 228232 3046 228482 3052
rect 228180 2994 228232 3000
rect 227352 2916 227404 2922
rect 227352 2858 227404 2864
rect 227536 2916 227588 2922
rect 227536 2858 227588 2864
rect 226340 2848 226392 2854
rect 226340 2790 226392 2796
rect 226352 480 226380 2790
rect 227548 480 227576 2858
rect 228744 480 228772 3062
rect 229572 2990 229600 3060
rect 229836 3052 229888 3058
rect 229836 2994 229888 3000
rect 229560 2984 229612 2990
rect 229560 2926 229612 2932
rect 229848 480 229876 2994
rect 230676 2854 230704 3060
rect 231032 2984 231084 2990
rect 231032 2926 231084 2932
rect 230664 2848 230716 2854
rect 230664 2790 230716 2796
rect 231044 480 231072 2926
rect 231780 2922 231808 3060
rect 232608 3046 232898 3062
rect 233712 3058 234002 3074
rect 233700 3052 234002 3058
rect 233752 3046 234002 3052
rect 234620 3052 234672 3058
rect 233700 2994 233752 3000
rect 234620 2994 234672 3000
rect 231768 2916 231820 2922
rect 231768 2858 231820 2864
rect 232228 2916 232280 2922
rect 232228 2858 232280 2864
rect 232240 480 232268 2858
rect 233424 2848 233476 2854
rect 233424 2790 233476 2796
rect 233436 480 233464 2790
rect 234632 480 234660 2994
rect 235092 2990 235120 3060
rect 235080 2984 235132 2990
rect 235080 2926 235132 2932
rect 235816 2984 235868 2990
rect 235816 2926 235868 2932
rect 235828 480 235856 2926
rect 236196 2922 236224 3060
rect 236184 2916 236236 2922
rect 236184 2858 236236 2864
rect 237012 2916 237064 2922
rect 237012 2858 237064 2864
rect 237024 480 237052 2858
rect 237300 2854 237328 3060
rect 238128 3058 238418 3074
rect 239312 3062 239364 3068
rect 242532 3120 242584 3126
rect 543464 3120 543516 3126
rect 242584 3068 242834 3074
rect 242532 3062 242834 3068
rect 238116 3052 238418 3058
rect 238168 3046 238418 3052
rect 238116 2994 238168 3000
rect 237288 2848 237340 2854
rect 237288 2790 237340 2796
rect 238116 2848 238168 2854
rect 238116 2790 238168 2796
rect 238128 480 238156 2790
rect 239324 480 239352 3062
rect 239508 2990 239536 3060
rect 240508 3052 240560 3058
rect 240508 2994 240560 3000
rect 239496 2984 239548 2990
rect 239496 2926 239548 2932
rect 240520 480 240548 2994
rect 240612 2922 240640 3060
rect 240600 2916 240652 2922
rect 240600 2858 240652 2864
rect 241716 2854 241744 3060
rect 242544 3046 242834 3062
rect 243648 3058 243938 3074
rect 243636 3052 243938 3058
rect 243688 3046 243938 3052
rect 243636 2994 243688 3000
rect 245028 2990 245056 3060
rect 245200 3052 245252 3058
rect 245200 2994 245252 3000
rect 242072 2984 242124 2990
rect 242072 2926 242124 2932
rect 245016 2984 245068 2990
rect 245016 2926 245068 2932
rect 241704 2848 241756 2854
rect 241704 2790 241756 2796
rect 222722 326 223160 354
rect 222722 -960 222834 326
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 354 241786 480
rect 242084 354 242112 2926
rect 244096 2916 244148 2922
rect 244096 2858 244148 2864
rect 242900 2848 242952 2854
rect 242900 2790 242952 2796
rect 242912 480 242940 2790
rect 244108 480 244136 2858
rect 245212 480 245240 2994
rect 246132 2854 246160 3060
rect 247236 2922 247264 3060
rect 248064 3058 248354 3074
rect 248052 3052 248354 3058
rect 248104 3046 248354 3052
rect 248788 3052 248840 3058
rect 248052 2994 248104 3000
rect 248788 2994 248840 3000
rect 247592 2984 247644 2990
rect 247592 2926 247644 2932
rect 247224 2916 247276 2922
rect 247224 2858 247276 2864
rect 246120 2848 246172 2854
rect 246120 2790 246172 2796
rect 246396 2848 246448 2854
rect 246396 2790 246448 2796
rect 246408 480 246436 2790
rect 247604 480 247632 2926
rect 248800 480 248828 2994
rect 249444 2854 249472 3060
rect 250548 2990 250576 3060
rect 251376 3058 251666 3074
rect 251364 3052 251666 3058
rect 251416 3046 251666 3052
rect 251364 2994 251416 3000
rect 250536 2984 250588 2990
rect 250536 2926 250588 2932
rect 252756 2922 252784 3060
rect 253480 2984 253532 2990
rect 253480 2926 253532 2932
rect 249984 2916 250036 2922
rect 249984 2858 250036 2864
rect 252744 2916 252796 2922
rect 252744 2858 252796 2864
rect 249432 2848 249484 2854
rect 249432 2790 249484 2796
rect 249996 480 250024 2858
rect 252376 2848 252428 2854
rect 252376 2790 252428 2796
rect 251180 808 251232 814
rect 251180 750 251232 756
rect 251192 480 251220 750
rect 252388 480 252416 2790
rect 253492 480 253520 2926
rect 253860 814 253888 3060
rect 254676 2916 254728 2922
rect 254676 2858 254728 2864
rect 253848 808 253900 814
rect 253848 750 253900 756
rect 254688 480 254716 2858
rect 254964 2854 254992 3060
rect 256068 2990 256096 3060
rect 256056 2984 256108 2990
rect 256056 2926 256108 2932
rect 257172 2922 257200 3060
rect 257160 2916 257212 2922
rect 257160 2858 257212 2864
rect 258276 2854 258304 3060
rect 254952 2848 255004 2854
rect 254952 2790 255004 2796
rect 255872 2848 255924 2854
rect 255872 2790 255924 2796
rect 258264 2848 258316 2854
rect 258264 2790 258316 2796
rect 255884 480 255912 2790
rect 259380 1358 259408 3060
rect 257068 1352 257120 1358
rect 257068 1294 257120 1300
rect 259368 1352 259420 1358
rect 259368 1294 259420 1300
rect 259460 1352 259512 1358
rect 259460 1294 259512 1300
rect 257080 480 257108 1294
rect 258264 1284 258316 1290
rect 258264 1226 258316 1232
rect 258276 480 258304 1226
rect 259472 480 259500 1294
rect 260484 1290 260512 3060
rect 260656 2848 260708 2854
rect 260656 2790 260708 2796
rect 260472 1284 260524 1290
rect 260472 1226 260524 1232
rect 260668 480 260696 2790
rect 261588 1358 261616 3060
rect 261760 2916 261812 2922
rect 261760 2858 261812 2864
rect 261576 1352 261628 1358
rect 261576 1294 261628 1300
rect 261772 480 261800 2858
rect 262692 2854 262720 3060
rect 263796 2922 263824 3060
rect 263784 2916 263836 2922
rect 263784 2858 263836 2864
rect 262680 2848 262732 2854
rect 262680 2790 262732 2796
rect 264900 1358 264928 3060
rect 262956 1352 263008 1358
rect 262956 1294 263008 1300
rect 264888 1352 264940 1358
rect 264888 1294 264940 1300
rect 265348 1352 265400 1358
rect 265348 1294 265400 1300
rect 262968 480 262996 1294
rect 264152 1284 264204 1290
rect 264152 1226 264204 1232
rect 264164 480 264192 1226
rect 265360 480 265388 1294
rect 266004 1290 266032 3060
rect 267108 1358 267136 3060
rect 267096 1352 267148 1358
rect 267096 1294 267148 1300
rect 267740 1352 267792 1358
rect 267740 1294 267792 1300
rect 265992 1284 266044 1290
rect 265992 1226 266044 1232
rect 266544 1284 266596 1290
rect 266544 1226 266596 1232
rect 266556 480 266584 1226
rect 267752 480 267780 1294
rect 268212 1290 268240 3060
rect 269316 1358 269344 3060
rect 269304 1352 269356 1358
rect 269304 1294 269356 1300
rect 268200 1284 268252 1290
rect 268200 1226 268252 1232
rect 270040 1284 270092 1290
rect 270040 1226 270092 1232
rect 268844 1216 268896 1222
rect 268844 1158 268896 1164
rect 268856 480 268884 1158
rect 270052 480 270080 1226
rect 270420 1222 270448 3060
rect 271236 1352 271288 1358
rect 271236 1294 271288 1300
rect 270408 1216 270460 1222
rect 270408 1158 270460 1164
rect 271248 480 271276 1294
rect 271524 1290 271552 3060
rect 272628 1358 272656 3060
rect 272616 1352 272668 1358
rect 272616 1294 272668 1300
rect 273628 1352 273680 1358
rect 273628 1294 273680 1300
rect 271512 1284 271564 1290
rect 271512 1226 271564 1232
rect 272432 1284 272484 1290
rect 272432 1226 272484 1232
rect 272444 480 272472 1226
rect 273640 480 273668 1294
rect 273732 1290 273760 3060
rect 274836 1358 274864 3060
rect 275296 3046 275954 3074
rect 276124 3046 277058 3074
rect 274824 1352 274876 1358
rect 274824 1294 274876 1300
rect 273720 1284 273772 1290
rect 273720 1226 273772 1232
rect 241674 326 242112 354
rect 241674 -960 241786 326
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 354 274906 480
rect 275296 354 275324 3046
rect 276124 1578 276152 3046
rect 276032 1550 276152 1578
rect 276032 480 276060 1550
rect 278148 1358 278176 3060
rect 278792 3046 279266 3074
rect 277124 1352 277176 1358
rect 277124 1294 277176 1300
rect 278136 1352 278188 1358
rect 278136 1294 278188 1300
rect 277136 480 277164 1294
rect 274794 326 275324 354
rect 274794 -960 274906 326
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 354 278402 480
rect 278792 354 278820 3046
rect 280356 1358 280384 3060
rect 281184 3046 281474 3074
rect 281920 3046 282578 3074
rect 283392 3046 283682 3074
rect 284312 3046 284786 3074
rect 285416 3046 285890 3074
rect 279516 1352 279568 1358
rect 279516 1294 279568 1300
rect 280344 1352 280396 1358
rect 280344 1294 280396 1300
rect 279528 480 279556 1294
rect 278290 326 278820 354
rect 278290 -960 278402 326
rect 279486 -960 279598 480
rect 280682 354 280794 480
rect 281184 354 281212 3046
rect 281920 480 281948 3046
rect 280682 326 281212 354
rect 280682 -960 280794 326
rect 281878 -960 281990 480
rect 283074 354 283186 480
rect 283392 354 283420 3046
rect 284312 480 284340 3046
rect 285416 480 285444 3046
rect 283074 326 283420 354
rect 283074 -960 283186 326
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 354 286682 480
rect 286980 354 287008 3060
rect 287808 3046 288098 3074
rect 287808 480 287836 3046
rect 286570 326 287008 354
rect 286570 -960 286682 326
rect 287766 -960 287878 480
rect 288962 354 289074 480
rect 289188 354 289216 3060
rect 290200 3046 290306 3074
rect 290200 480 290228 3046
rect 291396 480 291424 3060
rect 292592 480 292620 3060
rect 293696 480 293724 3060
rect 294814 3046 294920 3074
rect 294892 480 294920 3046
rect 288962 326 289216 354
rect 288962 -960 289074 326
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 295904 354 295932 3060
rect 297022 3046 297312 3074
rect 297284 480 297312 3046
rect 296046 354 296158 480
rect 295904 326 296158 354
rect 296046 -960 296158 326
rect 297242 -960 297354 480
rect 298112 354 298140 3060
rect 299230 3046 299704 3074
rect 300334 3046 300808 3074
rect 301438 3046 301728 3074
rect 302542 3046 303200 3074
rect 303646 3046 303936 3074
rect 299676 480 299704 3046
rect 300780 480 300808 3046
rect 298438 354 298550 480
rect 298112 326 298550 354
rect 298438 -960 298550 326
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301700 354 301728 3046
rect 303172 480 303200 3046
rect 301934 354 302046 480
rect 301700 326 302046 354
rect 301934 -960 302046 326
rect 303130 -960 303242 480
rect 303908 354 303936 3046
rect 304736 2854 304764 3060
rect 305854 3046 306328 3074
rect 304724 2848 304776 2854
rect 304724 2790 304776 2796
rect 305552 2848 305604 2854
rect 305552 2790 305604 2796
rect 305564 480 305592 2790
rect 304326 354 304438 480
rect 303908 326 304438 354
rect 304326 -960 304438 326
rect 305522 -960 305634 480
rect 306300 354 306328 3046
rect 306944 2854 306972 3060
rect 308062 3046 308996 3074
rect 306932 2848 306984 2854
rect 306932 2790 306984 2796
rect 307944 2848 307996 2854
rect 307944 2790 307996 2796
rect 307956 480 307984 2790
rect 308968 1578 308996 3046
rect 309152 2854 309180 3060
rect 310256 2990 310284 3060
rect 310244 2984 310296 2990
rect 310244 2926 310296 2932
rect 311360 2854 311388 3060
rect 311440 2984 311492 2990
rect 311440 2926 311492 2932
rect 309140 2848 309192 2854
rect 309140 2790 309192 2796
rect 310244 2848 310296 2854
rect 310244 2790 310296 2796
rect 311348 2848 311400 2854
rect 311348 2790 311400 2796
rect 308968 1550 309088 1578
rect 309060 480 309088 1550
rect 310256 480 310284 2790
rect 311452 480 311480 2926
rect 312464 2922 312492 3060
rect 312452 2916 312504 2922
rect 312452 2858 312504 2864
rect 313568 2854 313596 3060
rect 314580 2922 314608 3060
rect 313832 2916 313884 2922
rect 313832 2858 313884 2864
rect 314568 2916 314620 2922
rect 314568 2858 314620 2864
rect 312636 2848 312688 2854
rect 312636 2790 312688 2796
rect 313556 2848 313608 2854
rect 313556 2790 313608 2796
rect 312648 480 312676 2790
rect 313844 480 313872 2858
rect 315776 2854 315804 3060
rect 316880 2922 316908 3060
rect 316224 2916 316276 2922
rect 316224 2858 316276 2864
rect 316868 2916 316920 2922
rect 316868 2858 316920 2864
rect 315028 2848 315080 2854
rect 315028 2790 315080 2796
rect 315764 2848 315816 2854
rect 315764 2790 315816 2796
rect 315040 480 315068 2790
rect 316236 480 316264 2858
rect 317984 2854 318012 3060
rect 319088 2922 319116 3060
rect 318524 2916 318576 2922
rect 318524 2858 318576 2864
rect 319076 2916 319128 2922
rect 319076 2858 319128 2864
rect 317328 2848 317380 2854
rect 317328 2790 317380 2796
rect 317972 2848 318024 2854
rect 317972 2790 318024 2796
rect 317340 480 317368 2790
rect 318536 480 318564 2858
rect 320100 2854 320128 3060
rect 321296 2922 321324 3060
rect 320916 2916 320968 2922
rect 320916 2858 320968 2864
rect 321284 2916 321336 2922
rect 321284 2858 321336 2864
rect 319720 2848 319772 2854
rect 319720 2790 319772 2796
rect 320088 2848 320140 2854
rect 320088 2790 320140 2796
rect 319732 480 319760 2790
rect 320928 480 320956 2858
rect 322400 2854 322428 3060
rect 323504 2922 323532 3060
rect 323308 2916 323360 2922
rect 323308 2858 323360 2864
rect 323492 2916 323544 2922
rect 323492 2858 323544 2864
rect 322112 2848 322164 2854
rect 322112 2790 322164 2796
rect 322388 2848 322440 2854
rect 322388 2790 322440 2796
rect 322124 480 322152 2790
rect 323320 480 323348 2858
rect 324608 2854 324636 3060
rect 325712 2990 325740 3060
rect 326830 3046 327028 3074
rect 325700 2984 325752 2990
rect 325700 2926 325752 2932
rect 325608 2916 325660 2922
rect 325608 2858 325660 2864
rect 324412 2848 324464 2854
rect 324412 2790 324464 2796
rect 324596 2848 324648 2854
rect 324596 2790 324648 2796
rect 324424 480 324452 2790
rect 325620 480 325648 2858
rect 327000 2854 327028 3046
rect 327920 2922 327948 3060
rect 329024 2990 329052 3060
rect 328000 2984 328052 2990
rect 328000 2926 328052 2932
rect 329012 2984 329064 2990
rect 329012 2926 329064 2932
rect 327908 2916 327960 2922
rect 327908 2858 327960 2864
rect 326804 2848 326856 2854
rect 326804 2790 326856 2796
rect 326988 2848 327040 2854
rect 326988 2790 327040 2796
rect 326816 480 326844 2790
rect 328012 480 328040 2926
rect 330128 2854 330156 3060
rect 331140 2922 331168 3060
rect 332336 2990 332364 3060
rect 333454 3058 333744 3074
rect 333454 3052 333756 3058
rect 333454 3046 333704 3052
rect 333704 2994 333756 3000
rect 331588 2984 331640 2990
rect 331588 2926 331640 2932
rect 332324 2984 332376 2990
rect 332324 2926 332376 2932
rect 330392 2916 330444 2922
rect 330392 2858 330444 2864
rect 331128 2916 331180 2922
rect 331128 2858 331180 2864
rect 329196 2848 329248 2854
rect 329196 2790 329248 2796
rect 330116 2848 330168 2854
rect 330116 2790 330168 2796
rect 329208 480 329236 2790
rect 330404 480 330432 2858
rect 331600 480 331628 2926
rect 334544 2922 334572 3060
rect 335084 2984 335136 2990
rect 335084 2926 335136 2932
rect 333888 2916 333940 2922
rect 333888 2858 333940 2864
rect 334532 2916 334584 2922
rect 334532 2858 334584 2864
rect 332692 2848 332744 2854
rect 332692 2790 332744 2796
rect 332704 480 332732 2790
rect 333900 480 333928 2858
rect 335096 480 335124 2926
rect 335648 2854 335676 3060
rect 336280 3052 336332 3058
rect 336280 2994 336332 3000
rect 335636 2848 335688 2854
rect 335636 2790 335688 2796
rect 336292 480 336320 2994
rect 336660 1358 336688 3060
rect 337476 2916 337528 2922
rect 337476 2858 337528 2864
rect 336648 1352 336700 1358
rect 336648 1294 336700 1300
rect 337488 480 337516 2858
rect 337856 882 337884 3060
rect 338960 2854 338988 3060
rect 340064 2922 340092 3060
rect 341168 2990 341196 3060
rect 341156 2984 341208 2990
rect 341156 2926 341208 2932
rect 340052 2916 340104 2922
rect 340052 2858 340104 2864
rect 338672 2848 338724 2854
rect 338672 2790 338724 2796
rect 338948 2848 339000 2854
rect 338948 2790 339000 2796
rect 342076 2848 342128 2854
rect 342076 2790 342128 2796
rect 337844 876 337896 882
rect 337844 818 337896 824
rect 338684 480 338712 2790
rect 339868 1352 339920 1358
rect 339868 1294 339920 1300
rect 339880 480 339908 1294
rect 342088 1170 342116 2790
rect 342180 1358 342208 3060
rect 342996 2916 343048 2922
rect 342996 2858 343048 2864
rect 342168 1352 342220 1358
rect 342168 1294 342220 1300
rect 342088 1142 342208 1170
rect 340972 876 341024 882
rect 340972 818 341024 824
rect 340984 480 341012 818
rect 342180 480 342208 1142
rect 306718 354 306830 480
rect 306300 326 306830 354
rect 306718 -960 306830 326
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343008 354 343036 2858
rect 343376 1290 343404 3060
rect 344494 3046 344784 3074
rect 344560 2984 344612 2990
rect 344560 2926 344612 2932
rect 343364 1284 343416 1290
rect 343364 1226 343416 1232
rect 344572 480 344600 2926
rect 343334 354 343446 480
rect 343008 326 343446 354
rect 343334 -960 343446 326
rect 344530 -960 344642 480
rect 344756 66 344784 3046
rect 345584 1018 345612 3060
rect 346688 2854 346716 3060
rect 346676 2848 346728 2854
rect 346676 2790 346728 2796
rect 345756 1352 345808 1358
rect 345756 1294 345808 1300
rect 345572 1012 345624 1018
rect 345572 954 345624 960
rect 345768 480 345796 1294
rect 346952 1284 347004 1290
rect 346952 1226 347004 1232
rect 346964 480 346992 1226
rect 347700 882 347728 3060
rect 348896 1358 348924 3060
rect 348884 1352 348936 1358
rect 348884 1294 348936 1300
rect 350000 1290 350028 3060
rect 350448 2848 350500 2854
rect 350448 2790 350500 2796
rect 349988 1284 350040 1290
rect 349988 1226 350040 1232
rect 349252 1012 349304 1018
rect 349252 954 349304 960
rect 347688 876 347740 882
rect 347688 818 347740 824
rect 349264 480 349292 954
rect 350460 480 350488 2790
rect 351104 1018 351132 3060
rect 352208 1154 352236 3060
rect 353220 2854 353248 3060
rect 353208 2848 353260 2854
rect 353208 2790 353260 2796
rect 352840 1352 352892 1358
rect 352840 1294 352892 1300
rect 352196 1148 352248 1154
rect 352196 1090 352248 1096
rect 351092 1012 351144 1018
rect 351092 954 351144 960
rect 351644 876 351696 882
rect 351644 818 351696 824
rect 351656 480 351684 818
rect 352852 480 352880 1294
rect 354036 1284 354088 1290
rect 354036 1226 354088 1232
rect 354048 480 354076 1226
rect 344744 60 344796 66
rect 344744 2 344796 8
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 82 348138 480
rect 348026 66 348280 82
rect 348026 60 348292 66
rect 348026 54 348240 60
rect 348026 -960 348138 54
rect 348240 2 348292 8
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 354416 270 354444 3060
rect 355520 1086 355548 3060
rect 356624 1358 356652 3060
rect 357532 2848 357584 2854
rect 357532 2790 357584 2796
rect 356612 1352 356664 1358
rect 356612 1294 356664 1300
rect 356336 1148 356388 1154
rect 356336 1090 356388 1096
rect 355508 1080 355560 1086
rect 355508 1022 355560 1028
rect 355232 1012 355284 1018
rect 355232 954 355284 960
rect 355244 480 355272 954
rect 356348 480 356376 1090
rect 357544 480 357572 2790
rect 357728 1290 357756 3060
rect 357716 1284 357768 1290
rect 357716 1226 357768 1232
rect 358740 950 358768 3060
rect 359936 1222 359964 3060
rect 359924 1216 359976 1222
rect 359924 1158 359976 1164
rect 361040 1154 361068 3060
rect 361120 1352 361172 1358
rect 361120 1294 361172 1300
rect 361028 1148 361080 1154
rect 361028 1090 361080 1096
rect 359924 1080 359976 1086
rect 359924 1022 359976 1028
rect 358728 944 358780 950
rect 358728 886 358780 892
rect 359936 480 359964 1022
rect 361132 480 361160 1294
rect 362144 1018 362172 3060
rect 362316 1284 362368 1290
rect 362316 1226 362368 1232
rect 362132 1012 362184 1018
rect 362132 954 362184 960
rect 362328 480 362356 1226
rect 354404 264 354456 270
rect 354404 206 354456 212
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 218 358810 480
rect 358912 264 358964 270
rect 358698 212 358912 218
rect 358698 206 358964 212
rect 358698 190 358952 206
rect 358698 -960 358810 190
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363248 66 363276 3060
rect 364260 1358 364288 3060
rect 364248 1352 364300 1358
rect 364248 1294 364300 1300
rect 365456 1290 365484 3060
rect 365444 1284 365496 1290
rect 365444 1226 365496 1232
rect 366560 1222 366588 3060
rect 364616 1216 364668 1222
rect 364616 1158 364668 1164
rect 366548 1216 366600 1222
rect 366548 1158 366600 1164
rect 363512 944 363564 950
rect 363512 886 363564 892
rect 363524 480 363552 886
rect 364628 480 364656 1158
rect 367664 1154 367692 3060
rect 365444 1148 365496 1154
rect 365444 1090 365496 1096
rect 367652 1148 367704 1154
rect 367652 1090 367704 1096
rect 363236 60 363288 66
rect 363236 2 363288 8
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365456 354 365484 1090
rect 367008 1012 367060 1018
rect 367008 954 367060 960
rect 367020 480 367048 954
rect 368768 882 368796 3060
rect 369400 1352 369452 1358
rect 369400 1294 369452 1300
rect 368756 876 368808 882
rect 368756 818 368808 824
rect 369412 480 369440 1294
rect 369780 1018 369808 3060
rect 370976 1290 371004 3060
rect 372094 3046 372384 3074
rect 372356 2854 372384 3046
rect 372344 2848 372396 2854
rect 372344 2790 372396 2796
rect 370228 1284 370280 1290
rect 370228 1226 370280 1232
rect 370964 1284 371016 1290
rect 370964 1226 371016 1232
rect 369768 1012 369820 1018
rect 369768 954 369820 960
rect 365782 354 365894 480
rect 365456 326 365894 354
rect 365782 -960 365894 326
rect 366978 -960 367090 480
rect 368174 82 368286 480
rect 367848 66 368286 82
rect 367836 60 368286 66
rect 367888 54 368286 60
rect 367836 2 367888 8
rect 368174 -960 368286 54
rect 369370 -960 369482 480
rect 370240 354 370268 1226
rect 371332 1216 371384 1222
rect 371332 1158 371384 1164
rect 370566 354 370678 480
rect 370240 326 370678 354
rect 371344 354 371372 1158
rect 372896 1148 372948 1154
rect 372896 1090 372948 1096
rect 372908 480 372936 1090
rect 373184 1086 373212 3060
rect 374288 1358 374316 3060
rect 374276 1352 374328 1358
rect 374276 1294 374328 1300
rect 375300 1154 375328 3060
rect 376116 1284 376168 1290
rect 376116 1226 376168 1232
rect 375288 1148 375340 1154
rect 375288 1090 375340 1096
rect 373172 1080 373224 1086
rect 373172 1022 373224 1028
rect 375288 1012 375340 1018
rect 375288 954 375340 960
rect 373908 876 373960 882
rect 373908 818 373960 824
rect 371670 354 371782 480
rect 371344 326 371782 354
rect 370566 -960 370678 326
rect 371670 -960 371782 326
rect 372866 -960 372978 480
rect 373920 354 373948 818
rect 375300 480 375328 954
rect 374062 354 374174 480
rect 373920 326 374174 354
rect 374062 -960 374174 326
rect 375258 -960 375370 480
rect 376128 354 376156 1226
rect 376496 1018 376524 3060
rect 377600 1290 377628 3060
rect 377680 2848 377732 2854
rect 377680 2790 377732 2796
rect 377588 1284 377640 1290
rect 377588 1226 377640 1232
rect 376484 1012 376536 1018
rect 376484 954 376536 960
rect 377692 480 377720 2790
rect 378704 1222 378732 3060
rect 379612 1352 379664 1358
rect 379612 1294 379664 1300
rect 378692 1216 378744 1222
rect 378692 1158 378744 1164
rect 378508 1080 378560 1086
rect 378508 1022 378560 1028
rect 376454 354 376566 480
rect 376128 326 376566 354
rect 376454 -960 376566 326
rect 377650 -960 377762 480
rect 378520 354 378548 1022
rect 378846 354 378958 480
rect 378520 326 378958 354
rect 379624 354 379652 1294
rect 379808 1154 379836 3060
rect 379796 1148 379848 1154
rect 379796 1090 379848 1096
rect 379950 354 380062 480
rect 379624 326 380062 354
rect 378846 -960 378958 326
rect 379950 -960 380062 326
rect 380820 270 380848 3060
rect 381176 1080 381228 1086
rect 381176 1022 381228 1028
rect 381188 480 381216 1022
rect 380808 264 380860 270
rect 380808 206 380860 212
rect 381146 -960 381258 480
rect 382016 474 382044 3060
rect 382372 1012 382424 1018
rect 382372 954 382424 960
rect 382384 480 382412 954
rect 382004 468 382056 474
rect 382004 410 382056 416
rect 382342 -960 382454 480
rect 383120 66 383148 3060
rect 384224 1358 384252 3060
rect 384212 1352 384264 1358
rect 384212 1294 384264 1300
rect 383568 1284 383620 1290
rect 383568 1226 383620 1232
rect 383580 480 383608 1226
rect 384396 1216 384448 1222
rect 384396 1158 384448 1164
rect 383108 60 383160 66
rect 383108 2 383160 8
rect 383538 -960 383650 480
rect 384408 354 384436 1158
rect 385328 1086 385356 3060
rect 386340 1154 386368 3060
rect 387536 1222 387564 3060
rect 388640 1290 388668 3060
rect 388628 1284 388680 1290
rect 388628 1226 388680 1232
rect 387524 1216 387576 1222
rect 387524 1158 387576 1164
rect 385960 1148 386012 1154
rect 385960 1090 386012 1096
rect 386328 1148 386380 1154
rect 386328 1090 386380 1096
rect 385316 1080 385368 1086
rect 385316 1022 385368 1028
rect 385972 480 386000 1090
rect 389744 610 389772 3060
rect 390652 1352 390704 1358
rect 390652 1294 390704 1300
rect 389732 604 389784 610
rect 389732 546 389784 552
rect 390664 480 390692 1294
rect 384734 354 384846 480
rect 384408 326 384846 354
rect 384734 -960 384846 326
rect 385930 -960 386042 480
rect 386788 264 386840 270
rect 387126 218 387238 480
rect 387892 468 387944 474
rect 387892 410 387944 416
rect 387904 354 387932 410
rect 388230 354 388342 480
rect 387904 326 388342 354
rect 386840 212 387238 218
rect 386788 206 387238 212
rect 386800 190 387238 206
rect 387126 -960 387238 190
rect 388230 -960 388342 326
rect 389426 82 389538 480
rect 389426 66 389680 82
rect 389426 60 389692 66
rect 389426 54 389640 60
rect 389426 -960 389538 54
rect 389640 2 389692 8
rect 390622 -960 390734 480
rect 390848 66 390876 3060
rect 391676 3046 391874 3074
rect 391676 270 391704 3046
rect 392676 1148 392728 1154
rect 392676 1090 392728 1096
rect 391848 1080 391900 1086
rect 391848 1022 391900 1028
rect 391860 480 391888 1022
rect 391664 264 391716 270
rect 391664 206 391716 212
rect 390836 60 390888 66
rect 390836 2 390888 8
rect 391818 -960 391930 480
rect 392688 354 392716 1090
rect 393056 678 393084 3060
rect 394160 1086 394188 3060
rect 395264 1222 395292 3060
rect 396368 1358 396396 3060
rect 396356 1352 396408 1358
rect 396356 1294 396408 1300
rect 395344 1284 395396 1290
rect 395344 1226 395396 1232
rect 394240 1216 394292 1222
rect 394240 1158 394292 1164
rect 395252 1216 395304 1222
rect 395252 1158 395304 1164
rect 394148 1080 394200 1086
rect 394148 1022 394200 1028
rect 393044 672 393096 678
rect 393044 614 393096 620
rect 394252 480 394280 1158
rect 395356 480 395384 1226
rect 397380 1154 397408 3060
rect 397368 1148 397420 1154
rect 397368 1090 397420 1096
rect 396540 604 396592 610
rect 396540 546 396592 552
rect 396552 480 396580 546
rect 393014 354 393126 480
rect 392688 326 393126 354
rect 393014 -960 393126 326
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 82 397818 480
rect 398576 338 398604 3060
rect 398564 332 398616 338
rect 398564 274 398616 280
rect 398748 264 398800 270
rect 398902 218 399014 480
rect 398800 212 399014 218
rect 398748 206 399014 212
rect 398760 190 399014 206
rect 397706 66 397960 82
rect 397706 60 397972 66
rect 397706 54 397920 60
rect 397706 -960 397818 54
rect 397920 2 397972 8
rect 398902 -960 399014 190
rect 399680 134 399708 3060
rect 400784 678 400812 3060
rect 401324 1080 401376 1086
rect 401324 1022 401376 1028
rect 400128 672 400180 678
rect 400128 614 400180 620
rect 400772 672 400824 678
rect 400772 614 400824 620
rect 400140 480 400168 614
rect 401336 480 401364 1022
rect 401888 746 401916 3060
rect 402520 1216 402572 1222
rect 402520 1158 402572 1164
rect 401876 740 401928 746
rect 401876 682 401928 688
rect 402532 480 402560 1158
rect 399668 128 399720 134
rect 399668 70 399720 76
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 402900 66 402928 3060
rect 403624 1352 403676 1358
rect 403624 1294 403676 1300
rect 403636 480 403664 1294
rect 404096 1290 404124 3060
rect 404084 1284 404136 1290
rect 404084 1226 404136 1232
rect 404820 1148 404872 1154
rect 404820 1090 404872 1096
rect 404832 480 404860 1090
rect 402888 60 402940 66
rect 402888 2 402940 8
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405200 270 405228 3060
rect 406304 1358 406332 3060
rect 406292 1352 406344 1358
rect 406292 1294 406344 1300
rect 405986 354 406098 480
rect 405986 338 406240 354
rect 405986 332 406252 338
rect 405986 326 406200 332
rect 405188 264 405240 270
rect 405188 206 405240 212
rect 405986 -960 406098 326
rect 406200 274 406252 280
rect 407028 128 407080 134
rect 407182 82 407294 480
rect 407408 406 407436 3060
rect 408420 610 408448 3060
rect 409236 740 409288 746
rect 409236 682 409288 688
rect 408592 672 408644 678
rect 408592 614 408644 620
rect 408408 604 408460 610
rect 408408 546 408460 552
rect 407396 400 407448 406
rect 407396 342 407448 348
rect 407080 76 407294 82
rect 407028 70 407294 76
rect 407040 54 407294 70
rect 407182 -960 407294 54
rect 408378 218 408490 480
rect 408604 218 408632 614
rect 408378 190 408632 218
rect 409248 218 409276 682
rect 409616 678 409644 3060
rect 410734 3046 411024 3074
rect 411838 3046 412128 3074
rect 409604 672 409656 678
rect 409604 614 409656 620
rect 409574 218 409686 480
rect 409248 190 409686 218
rect 408378 -960 408490 190
rect 409574 -960 409686 190
rect 410770 82 410882 480
rect 410996 338 411024 3046
rect 411904 1284 411956 1290
rect 411904 1226 411956 1232
rect 411916 480 411944 1226
rect 410984 332 411036 338
rect 410984 274 411036 280
rect 410770 66 411024 82
rect 410770 60 411036 66
rect 410770 54 410984 60
rect 410770 -960 410882 54
rect 410984 2 411036 8
rect 411874 -960 411986 480
rect 412100 474 412128 3046
rect 412928 1222 412956 3060
rect 413940 1290 413968 3060
rect 414296 1352 414348 1358
rect 414296 1294 414348 1300
rect 413928 1284 413980 1290
rect 413928 1226 413980 1232
rect 412916 1216 412968 1222
rect 412916 1158 412968 1164
rect 414308 480 414336 1294
rect 415136 1086 415164 3060
rect 415124 1080 415176 1086
rect 415124 1022 415176 1028
rect 416240 950 416268 3060
rect 416228 944 416280 950
rect 416228 886 416280 892
rect 416688 604 416740 610
rect 416688 546 416740 552
rect 416700 480 416728 546
rect 412088 468 412140 474
rect 412088 410 412140 416
rect 412824 264 412876 270
rect 413070 218 413182 480
rect 412876 212 413182 218
rect 412824 206 413182 212
rect 412836 190 413182 206
rect 413070 -960 413182 190
rect 414266 -960 414378 480
rect 415308 400 415360 406
rect 415462 354 415574 480
rect 415360 348 415574 354
rect 415308 342 415574 348
rect 415320 326 415574 342
rect 415462 -960 415574 326
rect 416658 -960 416770 480
rect 417344 66 417372 3060
rect 417884 672 417936 678
rect 417884 614 417936 620
rect 417896 480 417924 614
rect 417332 60 417384 66
rect 417332 2 417384 8
rect 417854 -960 417966 480
rect 418448 202 418476 3060
rect 419460 1358 419488 3060
rect 419448 1352 419500 1358
rect 419448 1294 419500 1300
rect 420656 1154 420684 3060
rect 421760 1222 421788 3060
rect 422576 1284 422628 1290
rect 422576 1226 422628 1232
rect 421380 1216 421432 1222
rect 421380 1158 421432 1164
rect 421748 1216 421800 1222
rect 421748 1158 421800 1164
rect 420644 1148 420696 1154
rect 420644 1090 420696 1096
rect 421392 480 421420 1158
rect 422588 480 422616 1226
rect 422864 1018 422892 3060
rect 423404 1080 423456 1086
rect 423404 1022 423456 1028
rect 422852 1012 422904 1018
rect 422852 954 422904 960
rect 418958 354 419070 480
rect 418632 338 419070 354
rect 418620 332 419070 338
rect 418672 326 419070 332
rect 418620 274 418672 280
rect 418436 196 418488 202
rect 418436 138 418488 144
rect 418958 -960 419070 326
rect 420154 354 420266 480
rect 420368 468 420420 474
rect 420368 410 420420 416
rect 420380 354 420408 410
rect 420154 326 420408 354
rect 420154 -960 420266 326
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423416 354 423444 1022
rect 423742 354 423854 480
rect 423416 326 423854 354
rect 423742 -960 423854 326
rect 423968 134 423996 3060
rect 424980 1086 425008 3060
rect 426176 1290 426204 3060
rect 426164 1284 426216 1290
rect 426164 1226 426216 1232
rect 424968 1080 425020 1086
rect 424968 1022 425020 1028
rect 424968 944 425020 950
rect 424968 886 425020 892
rect 424980 480 425008 886
rect 427280 814 427308 3060
rect 428384 1358 428412 3060
rect 428280 1352 428332 1358
rect 428280 1294 428332 1300
rect 428372 1352 428424 1358
rect 428372 1294 428424 1300
rect 427268 808 427320 814
rect 427268 750 427320 756
rect 428292 762 428320 1294
rect 429292 1148 429344 1154
rect 429292 1090 429344 1096
rect 428292 734 428504 762
rect 428476 480 428504 734
rect 423956 128 424008 134
rect 423956 70 424008 76
rect 424938 -960 425050 480
rect 426134 82 426246 480
rect 427238 218 427350 480
rect 426912 202 427350 218
rect 426900 196 427350 202
rect 426952 190 427350 196
rect 426900 138 426952 144
rect 425808 66 426246 82
rect 425796 60 426246 66
rect 425848 54 426246 60
rect 425796 2 425848 8
rect 426134 -960 426246 54
rect 427238 -960 427350 190
rect 428434 -960 428546 480
rect 429304 354 429332 1090
rect 429488 746 429516 3060
rect 429476 740 429528 746
rect 429476 682 429528 688
rect 430500 542 430528 3060
rect 430856 1216 430908 1222
rect 430856 1158 430908 1164
rect 430488 536 430540 542
rect 429630 354 429742 480
rect 430488 478 430540 484
rect 430868 480 430896 1158
rect 431696 610 431724 3060
rect 432800 1018 432828 3060
rect 431868 1012 431920 1018
rect 431868 954 431920 960
rect 432788 1012 432840 1018
rect 432788 954 432840 960
rect 431684 604 431736 610
rect 431684 546 431736 552
rect 429304 326 429742 354
rect 429630 -960 429742 326
rect 430826 -960 430938 480
rect 431880 354 431908 954
rect 433904 950 433932 3060
rect 435008 1154 435036 3060
rect 436020 1358 436048 3060
rect 436008 1352 436060 1358
rect 436008 1294 436060 1300
rect 435180 1284 435232 1290
rect 435180 1226 435232 1232
rect 434996 1148 435048 1154
rect 434996 1090 435048 1096
rect 434076 1080 434128 1086
rect 434076 1022 434128 1028
rect 433892 944 433944 950
rect 433892 886 433944 892
rect 432022 354 432134 480
rect 431880 326 432134 354
rect 432022 -960 432134 326
rect 433218 82 433330 480
rect 434088 354 434116 1022
rect 434414 354 434526 480
rect 434088 326 434526 354
rect 435192 354 435220 1226
rect 436744 808 436796 814
rect 436744 750 436796 756
rect 436756 480 436784 750
rect 435518 354 435630 480
rect 435192 326 435630 354
rect 433432 128 433484 134
rect 433218 76 433432 82
rect 433218 70 433484 76
rect 433218 54 433472 70
rect 433218 -960 433330 54
rect 434414 -960 434526 326
rect 435518 -960 435630 326
rect 436714 -960 436826 480
rect 437216 474 437244 3060
rect 438320 1290 438348 3060
rect 437572 1284 437624 1290
rect 437572 1226 437624 1232
rect 438308 1284 438360 1290
rect 438308 1226 438360 1232
rect 437204 468 437256 474
rect 437204 410 437256 416
rect 437584 354 437612 1226
rect 439424 1222 439452 3060
rect 439412 1216 439464 1222
rect 439412 1158 439464 1164
rect 440528 746 440556 3060
rect 441540 1086 441568 3060
rect 441528 1080 441580 1086
rect 441528 1022 441580 1028
rect 442632 1012 442684 1018
rect 442632 954 442684 960
rect 439136 740 439188 746
rect 439136 682 439188 688
rect 440516 740 440568 746
rect 440516 682 440568 688
rect 439148 480 439176 682
rect 441528 672 441580 678
rect 441528 614 441580 620
rect 440332 604 440384 610
rect 440332 546 440384 552
rect 440344 480 440372 546
rect 441540 480 441568 614
rect 442644 480 442672 954
rect 442736 814 442764 3060
rect 443840 1358 443868 3060
rect 444958 3046 445248 3074
rect 443828 1352 443880 1358
rect 443828 1294 443880 1300
rect 443552 1216 443604 1222
rect 443552 1158 443604 1164
rect 443564 1018 443592 1158
rect 445220 1154 445248 3046
rect 445852 1284 445904 1290
rect 445852 1226 445904 1232
rect 445024 1148 445076 1154
rect 445024 1090 445076 1096
rect 445208 1148 445260 1154
rect 445208 1090 445260 1096
rect 443552 1012 443604 1018
rect 443552 954 443604 960
rect 443460 944 443512 950
rect 443460 886 443512 892
rect 442724 808 442776 814
rect 442724 750 442776 756
rect 437910 354 438022 480
rect 437584 326 438022 354
rect 437910 -960 438022 326
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443472 354 443500 886
rect 445036 480 445064 1090
rect 443798 354 443910 480
rect 443472 326 443910 354
rect 443798 -960 443910 326
rect 444994 -960 445106 480
rect 445864 354 445892 1226
rect 446048 950 446076 3060
rect 446036 944 446088 950
rect 446036 886 446088 892
rect 447060 610 447088 3060
rect 448256 882 448284 3060
rect 449360 1290 449388 3060
rect 449348 1284 449400 1290
rect 449348 1226 449400 1232
rect 450464 1222 450492 3060
rect 448612 1216 448664 1222
rect 448612 1158 448664 1164
rect 450452 1216 450504 1222
rect 450452 1158 450504 1164
rect 448244 876 448296 882
rect 448244 818 448296 824
rect 447048 604 447100 610
rect 447048 546 447100 552
rect 447244 598 447456 626
rect 446190 354 446302 480
rect 447244 474 447272 598
rect 447428 480 447456 598
rect 448624 480 448652 1158
rect 449808 1012 449860 1018
rect 449808 954 449860 960
rect 449820 480 449848 954
rect 451568 746 451596 3060
rect 451740 1080 451792 1086
rect 451740 1022 451792 1028
rect 450912 740 450964 746
rect 450912 682 450964 688
rect 451556 740 451608 746
rect 451556 682 451608 688
rect 450924 480 450952 682
rect 447232 468 447284 474
rect 447232 410 447284 416
rect 445864 326 446302 354
rect 446190 -960 446302 326
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 451752 354 451780 1022
rect 452078 354 452190 480
rect 451752 326 452190 354
rect 452078 -960 452190 326
rect 452580 134 452608 3060
rect 453304 808 453356 814
rect 453304 750 453356 756
rect 453316 480 453344 750
rect 452568 128 452620 134
rect 452568 70 452620 76
rect 453274 -960 453386 480
rect 453776 338 453804 3060
rect 454132 1352 454184 1358
rect 454132 1294 454184 1300
rect 454144 354 454172 1294
rect 454880 1290 454908 3060
rect 454868 1284 454920 1290
rect 454868 1226 454920 1232
rect 455696 1148 455748 1154
rect 455696 1090 455748 1096
rect 455708 480 455736 1090
rect 455984 1086 456012 3060
rect 457088 1358 457116 3060
rect 457916 3046 458114 3074
rect 459310 3046 459508 3074
rect 460414 3046 460612 3074
rect 456984 1352 457036 1358
rect 456984 1294 457036 1300
rect 457076 1352 457128 1358
rect 457076 1294 457128 1300
rect 455972 1080 456024 1086
rect 455972 1022 456024 1028
rect 456892 944 456944 950
rect 456892 886 456944 892
rect 456904 480 456932 886
rect 456996 678 457024 1294
rect 456984 672 457036 678
rect 456984 614 457036 620
rect 454470 354 454582 480
rect 453764 332 453816 338
rect 454144 326 454582 354
rect 453764 274 453816 280
rect 454470 -960 454582 326
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 457916 270 457944 3046
rect 459192 876 459244 882
rect 459192 818 459244 824
rect 458088 604 458140 610
rect 458088 546 458140 552
rect 458100 480 458128 546
rect 459204 480 459232 818
rect 459480 542 459508 3046
rect 460020 672 460072 678
rect 460020 614 460072 620
rect 459468 536 459520 542
rect 457904 264 457956 270
rect 457904 206 457956 212
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 459468 478 459520 484
rect 460032 354 460060 614
rect 460358 354 460470 480
rect 460584 406 460612 3046
rect 461504 610 461532 3060
rect 462608 1290 462636 3060
rect 462596 1284 462648 1290
rect 462596 1226 462648 1232
rect 461584 1148 461636 1154
rect 461584 1090 461636 1096
rect 461492 604 461544 610
rect 461492 546 461544 552
rect 461596 480 461624 1090
rect 462412 808 462464 814
rect 462412 750 462464 756
rect 460032 326 460470 354
rect 460572 400 460624 406
rect 460572 342 460624 348
rect 460358 -960 460470 326
rect 461554 -960 461666 480
rect 462424 354 462452 750
rect 462750 354 462862 480
rect 462424 326 462862 354
rect 462750 -960 462862 326
rect 463620 66 463648 3060
rect 464816 678 464844 3060
rect 464804 672 464856 678
rect 464804 614 464856 620
rect 463946 82 464058 480
rect 465142 354 465254 480
rect 465000 338 465254 354
rect 464988 332 465254 338
rect 465040 326 465254 332
rect 464988 274 465040 280
rect 464160 128 464212 134
rect 463946 76 464160 82
rect 463946 70 464212 76
rect 463608 60 463660 66
rect 463608 2 463660 8
rect 463946 54 464200 70
rect 463946 -960 464058 54
rect 465142 -960 465254 326
rect 465828 202 465856 3060
rect 465908 1216 465960 1222
rect 465908 1158 465960 1164
rect 465920 354 465948 1158
rect 466246 354 466358 480
rect 465920 326 466358 354
rect 465816 196 465868 202
rect 465816 138 465868 144
rect 466246 -960 466358 326
rect 467024 134 467052 3060
rect 467472 1080 467524 1086
rect 467472 1022 467524 1028
rect 467484 480 467512 1022
rect 468128 746 468156 3060
rect 468300 1352 468352 1358
rect 468300 1294 468352 1300
rect 468116 740 468168 746
rect 468116 682 468168 688
rect 467012 128 467064 134
rect 467012 70 467064 76
rect 467442 -960 467554 480
rect 468312 354 468340 1294
rect 469140 1154 469168 3060
rect 469128 1148 469180 1154
rect 469128 1090 469180 1096
rect 468638 354 468750 480
rect 468312 326 468750 354
rect 468638 -960 468750 326
rect 469834 218 469946 480
rect 470336 474 470364 3060
rect 470784 536 470836 542
rect 470784 478 470836 484
rect 470324 468 470376 474
rect 470324 410 470376 416
rect 470796 354 470824 478
rect 471030 354 471142 480
rect 470796 326 471142 354
rect 471440 338 471468 3060
rect 472226 354 472338 480
rect 472440 400 472492 406
rect 472226 348 472440 354
rect 472226 342 472492 348
rect 470048 264 470100 270
rect 469834 212 470048 218
rect 469834 206 470100 212
rect 469834 190 470088 206
rect 469834 -960 469946 190
rect 471030 -960 471142 326
rect 471428 332 471480 338
rect 471428 274 471480 280
rect 472226 326 472480 342
rect 472226 -960 472338 326
rect 472544 270 472572 3060
rect 473452 604 473504 610
rect 473452 546 473504 552
rect 473464 480 473492 546
rect 473648 542 473676 3060
rect 474188 1284 474240 1290
rect 474188 1226 474240 1232
rect 473636 536 473688 542
rect 472532 264 472584 270
rect 472532 206 472584 212
rect 473422 -960 473534 480
rect 473636 478 473688 484
rect 474200 354 474228 1226
rect 474660 1086 474688 3060
rect 475856 1222 475884 3060
rect 476974 3046 477264 3074
rect 478078 3046 478368 3074
rect 475844 1216 475896 1222
rect 475844 1158 475896 1164
rect 474648 1080 474700 1086
rect 474648 1022 474700 1028
rect 476948 672 477000 678
rect 476948 614 477000 620
rect 476960 480 476988 614
rect 474526 354 474638 480
rect 474200 326 474638 354
rect 474526 -960 474638 326
rect 475722 82 475834 480
rect 475722 66 475976 82
rect 475722 60 475988 66
rect 475722 54 475936 60
rect 475722 -960 475834 54
rect 475936 2 475988 8
rect 476918 -960 477030 480
rect 477236 66 477264 3046
rect 478114 218 478226 480
rect 478340 406 478368 3046
rect 478328 400 478380 406
rect 478328 342 478380 348
rect 478114 202 478368 218
rect 479168 202 479196 3060
rect 480180 1290 480208 3060
rect 481376 1358 481404 3060
rect 481364 1352 481416 1358
rect 481364 1294 481416 1300
rect 480168 1284 480220 1290
rect 480168 1226 480220 1232
rect 481364 1148 481416 1154
rect 481364 1090 481416 1096
rect 480536 740 480588 746
rect 480536 682 480588 688
rect 480548 480 480576 682
rect 478114 196 478380 202
rect 478114 190 478328 196
rect 477224 60 477276 66
rect 477224 2 477276 8
rect 478114 -960 478226 190
rect 478328 138 478380 144
rect 479156 196 479208 202
rect 479156 138 479208 144
rect 478972 128 479024 134
rect 479310 82 479422 480
rect 479024 76 479422 82
rect 478972 70 479422 76
rect 478984 54 479422 70
rect 479310 -960 479422 54
rect 480506 -960 480618 480
rect 481376 354 481404 1090
rect 482480 746 482508 3060
rect 483584 814 483612 3060
rect 483572 808 483624 814
rect 483572 750 483624 756
rect 482468 740 482520 746
rect 482468 682 482520 688
rect 481702 354 481814 480
rect 482468 468 482520 474
rect 482468 410 482520 416
rect 481376 326 481814 354
rect 482480 354 482508 410
rect 482806 354 482918 480
rect 482480 326 482918 354
rect 481702 -960 481814 326
rect 482806 -960 482918 326
rect 484002 354 484114 480
rect 484688 474 484716 3060
rect 485700 882 485728 3060
rect 485688 876 485740 882
rect 485688 818 485740 824
rect 486896 678 486924 3060
rect 488000 1154 488028 3060
rect 488816 1216 488868 1222
rect 488816 1158 488868 1164
rect 487988 1148 488040 1154
rect 487988 1090 488040 1096
rect 487252 1080 487304 1086
rect 487252 1022 487304 1028
rect 486884 672 486936 678
rect 486884 614 486936 620
rect 486424 604 486476 610
rect 486424 546 486476 552
rect 486436 480 486464 546
rect 484676 468 484728 474
rect 484676 410 484728 416
rect 484002 338 484256 354
rect 484002 332 484268 338
rect 484002 326 484216 332
rect 484002 -960 484114 326
rect 484216 274 484268 280
rect 484860 264 484912 270
rect 485198 218 485310 480
rect 484912 212 485310 218
rect 484860 206 485310 212
rect 484872 190 485310 206
rect 485198 -960 485310 190
rect 486394 -960 486506 480
rect 487264 354 487292 1022
rect 488828 480 488856 1158
rect 489104 1018 489132 3060
rect 489092 1012 489144 1018
rect 489092 954 489144 960
rect 487590 354 487702 480
rect 487264 326 487702 354
rect 487590 -960 487702 326
rect 488786 -960 488898 480
rect 489890 82 490002 480
rect 490208 474 490236 3060
rect 491220 626 491248 3060
rect 492430 3046 492628 3074
rect 491220 598 491340 626
rect 490196 468 490248 474
rect 490196 410 490248 416
rect 490748 400 490800 406
rect 491086 354 491198 480
rect 490800 348 491198 354
rect 490748 342 491198 348
rect 490760 326 491198 342
rect 489890 66 490144 82
rect 489890 60 490156 66
rect 489890 54 490104 60
rect 489890 -960 490002 54
rect 490104 2 490156 8
rect 491086 -960 491198 326
rect 491312 134 491340 598
rect 492282 218 492394 480
rect 492282 202 492536 218
rect 492600 202 492628 3046
rect 493520 1290 493548 3060
rect 493140 1284 493192 1290
rect 493140 1226 493192 1232
rect 493508 1284 493560 1290
rect 493508 1226 493560 1232
rect 493152 354 493180 1226
rect 494624 950 494652 3060
rect 495728 1358 495756 3060
rect 494704 1352 494756 1358
rect 494704 1294 494756 1300
rect 495716 1352 495768 1358
rect 495716 1294 495768 1300
rect 494612 944 494664 950
rect 494612 886 494664 892
rect 494716 480 494744 1294
rect 495532 740 495584 746
rect 495532 682 495584 688
rect 493478 354 493590 480
rect 493152 326 493590 354
rect 492282 196 492548 202
rect 492282 190 492496 196
rect 491300 128 491352 134
rect 491300 70 491352 76
rect 492282 -960 492394 190
rect 492496 138 492548 144
rect 492588 196 492640 202
rect 492588 138 492640 144
rect 493478 -960 493590 326
rect 494674 -960 494786 480
rect 495544 354 495572 682
rect 495870 354 495982 480
rect 495544 326 495982 354
rect 495870 -960 495982 326
rect 496740 66 496768 3060
rect 497096 808 497148 814
rect 497096 750 497148 756
rect 497108 480 497136 750
rect 496728 60 496780 66
rect 496728 2 496780 8
rect 497066 -960 497178 480
rect 497936 406 497964 3060
rect 498936 876 498988 882
rect 498936 818 498988 824
rect 498200 604 498252 610
rect 498200 546 498252 552
rect 498212 480 498240 546
rect 497924 400 497976 406
rect 497924 342 497976 348
rect 498170 -960 498282 480
rect 498948 354 498976 818
rect 499040 814 499068 3060
rect 499028 808 499080 814
rect 499028 750 499080 756
rect 499366 354 499478 480
rect 500144 474 500172 3060
rect 501248 1222 501276 3060
rect 501236 1216 501288 1222
rect 501236 1158 501288 1164
rect 501420 1148 501472 1154
rect 501420 1090 501472 1096
rect 500592 672 500644 678
rect 500592 614 500644 620
rect 500604 480 500632 614
rect 500132 468 500184 474
rect 500132 410 500184 416
rect 498948 326 499478 354
rect 499366 -960 499478 326
rect 500562 -960 500674 480
rect 501432 354 501460 1090
rect 502260 746 502288 3060
rect 502984 1012 503036 1018
rect 502984 954 503036 960
rect 502248 740 502300 746
rect 502248 682 502300 688
rect 502996 480 503024 954
rect 503456 678 503484 3060
rect 503444 672 503496 678
rect 503444 614 503496 620
rect 503812 604 503864 610
rect 503812 546 503864 552
rect 501758 354 501870 480
rect 501432 326 501870 354
rect 501758 -960 501870 326
rect 502954 -960 503066 480
rect 503824 354 503852 546
rect 504150 354 504262 480
rect 504560 406 504588 3060
rect 503824 326 504262 354
rect 504548 400 504600 406
rect 504548 342 504600 348
rect 504150 -960 504262 326
rect 505346 82 505458 480
rect 505664 338 505692 3060
rect 506768 1154 506796 3060
rect 507780 1290 507808 3060
rect 507308 1284 507360 1290
rect 507308 1226 507360 1232
rect 507768 1284 507820 1290
rect 507768 1226 507820 1232
rect 506756 1148 506808 1154
rect 506756 1090 506808 1096
rect 505652 332 505704 338
rect 505652 274 505704 280
rect 506450 218 506562 480
rect 507320 354 507348 1226
rect 508872 944 508924 950
rect 508872 886 508924 892
rect 508884 480 508912 886
rect 508976 610 509004 3060
rect 510080 1358 510108 3060
rect 511198 3046 511488 3074
rect 512302 3046 512684 3074
rect 509700 1352 509752 1358
rect 509700 1294 509752 1300
rect 510068 1352 510120 1358
rect 510068 1294 510120 1300
rect 508964 604 509016 610
rect 508964 546 509016 552
rect 507646 354 507758 480
rect 507320 326 507758 354
rect 506450 202 506704 218
rect 506450 196 506716 202
rect 506450 190 506664 196
rect 505560 128 505612 134
rect 505346 76 505560 82
rect 505346 70 505612 76
rect 505346 54 505600 70
rect 505346 -960 505458 54
rect 506450 -960 506562 190
rect 506664 138 506716 144
rect 507646 -960 507758 326
rect 508842 -960 508954 480
rect 509712 354 509740 1294
rect 510038 354 510150 480
rect 509712 326 510150 354
rect 510038 -960 510150 326
rect 511234 82 511346 480
rect 511460 270 511488 3046
rect 512092 536 512144 542
rect 512092 478 512144 484
rect 512104 354 512132 478
rect 512430 354 512542 480
rect 512104 326 512542 354
rect 511448 264 511500 270
rect 511448 206 511500 212
rect 511234 66 511488 82
rect 511234 60 511500 66
rect 511234 54 511448 60
rect 511234 -960 511346 54
rect 511448 2 511500 8
rect 512430 -960 512542 326
rect 512656 202 512684 3046
rect 513300 2990 513328 3060
rect 513288 2984 513340 2990
rect 513288 2926 513340 2932
rect 513564 808 513616 814
rect 513564 750 513616 756
rect 513576 480 513604 750
rect 512644 196 512696 202
rect 512644 138 512696 144
rect 513534 -960 513646 480
rect 514496 134 514524 3060
rect 515496 1216 515548 1222
rect 515496 1158 515548 1164
rect 514730 354 514842 480
rect 514944 468 514996 474
rect 514944 410 514996 416
rect 514956 354 514984 410
rect 514730 326 514984 354
rect 515508 354 515536 1158
rect 515600 950 515628 3060
rect 516704 1222 516732 3060
rect 517520 2916 517572 2922
rect 517520 2858 517572 2864
rect 517532 1290 517560 2858
rect 517612 2848 517664 2854
rect 517612 2790 517664 2796
rect 517520 1284 517572 1290
rect 517520 1226 517572 1232
rect 516692 1216 516744 1222
rect 516692 1158 516744 1164
rect 517624 1154 517652 2790
rect 517612 1148 517664 1154
rect 517612 1090 517664 1096
rect 515588 944 515640 950
rect 515588 886 515640 892
rect 517152 740 517204 746
rect 517152 682 517204 688
rect 517164 480 517192 682
rect 517808 542 517836 3060
rect 518820 1086 518848 3060
rect 518808 1080 518860 1086
rect 518808 1022 518860 1028
rect 520016 1018 520044 3060
rect 520004 1012 520056 1018
rect 520004 954 520056 960
rect 521120 746 521148 3060
rect 521844 2848 521896 2854
rect 521844 2790 521896 2796
rect 521108 740 521160 746
rect 521108 682 521160 688
rect 518348 672 518400 678
rect 518348 614 518400 620
rect 517796 536 517848 542
rect 515926 354 516038 480
rect 515508 326 516038 354
rect 514484 128 514536 134
rect 514484 70 514536 76
rect 514730 -960 514842 326
rect 515926 -960 516038 326
rect 517122 -960 517234 480
rect 517796 478 517848 484
rect 518360 480 518388 614
rect 521856 480 521884 2790
rect 522224 1154 522252 3060
rect 523040 2916 523092 2922
rect 523040 2858 523092 2864
rect 522212 1148 522264 1154
rect 522212 1090 522264 1096
rect 523052 480 523080 2858
rect 523328 678 523356 3060
rect 524340 678 524368 3060
rect 525550 3046 525748 3074
rect 526654 3046 526944 3074
rect 525432 1352 525484 1358
rect 525432 1294 525484 1300
rect 523316 672 523368 678
rect 523316 614 523368 620
rect 524328 672 524380 678
rect 524328 614 524380 620
rect 523868 604 523920 610
rect 523868 546 523920 552
rect 518318 -960 518430 480
rect 519514 354 519626 480
rect 519728 400 519780 406
rect 519514 348 519728 354
rect 520710 354 520822 480
rect 519514 342 519780 348
rect 519514 326 519768 342
rect 520384 338 520822 354
rect 520372 332 520822 338
rect 519514 -960 519626 326
rect 520424 326 520822 332
rect 520372 274 520424 280
rect 520710 -960 520822 326
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 523880 354 523908 546
rect 525444 480 525472 1294
rect 524206 354 524318 480
rect 523880 326 524318 354
rect 524206 -960 524318 326
rect 525402 -960 525514 480
rect 525720 474 525748 3046
rect 525800 2916 525852 2922
rect 525800 2858 525852 2864
rect 525812 950 525840 2858
rect 525800 944 525852 950
rect 525800 886 525852 892
rect 525708 468 525760 474
rect 525708 410 525760 416
rect 526260 264 526312 270
rect 526598 218 526710 480
rect 526312 212 526710 218
rect 526260 206 526710 212
rect 526272 190 526710 206
rect 526598 -960 526710 190
rect 526916 66 526944 3046
rect 527744 882 527772 3060
rect 527732 876 527784 882
rect 527732 818 527784 824
rect 528848 814 528876 3060
rect 529966 3058 530072 3074
rect 529966 3052 530084 3058
rect 529966 3046 530032 3052
rect 530032 2994 530084 3000
rect 529020 2984 529072 2990
rect 529020 2926 529072 2932
rect 528836 808 528888 814
rect 528836 750 528888 756
rect 529032 480 529060 2926
rect 527794 218 527906 480
rect 527794 202 528048 218
rect 527794 196 528060 202
rect 527794 190 528008 196
rect 526904 60 526956 66
rect 526904 2 526956 8
rect 527794 -960 527906 190
rect 528008 138 528060 144
rect 528990 -960 529102 480
rect 529940 128 529992 134
rect 530094 82 530206 480
rect 531056 338 531084 3060
rect 531320 2916 531372 2922
rect 531320 2858 531372 2864
rect 531332 480 531360 2858
rect 532056 1216 532108 1222
rect 532056 1158 532108 1164
rect 531044 332 531096 338
rect 531044 274 531096 280
rect 529992 76 530206 82
rect 529940 70 530206 76
rect 529952 54 530206 70
rect 530094 -960 530206 54
rect 531290 -960 531402 480
rect 532068 354 532096 1158
rect 532160 950 532188 3060
rect 533278 3046 533844 3074
rect 543214 3068 543464 3074
rect 560484 3120 560536 3126
rect 543214 3062 543516 3068
rect 532148 944 532200 950
rect 532148 886 532200 892
rect 533252 672 533304 678
rect 533252 614 533304 620
rect 532486 354 532598 480
rect 533264 406 533292 614
rect 533816 610 533844 3046
rect 534368 1290 534396 3060
rect 534356 1284 534408 1290
rect 534356 1226 534408 1232
rect 534540 1080 534592 1086
rect 534540 1022 534592 1028
rect 533712 604 533764 610
rect 533712 546 533764 552
rect 533804 604 533856 610
rect 533804 546 533856 552
rect 533724 480 533752 546
rect 532068 326 532598 354
rect 533252 400 533304 406
rect 533252 342 533304 348
rect 532486 -960 532598 326
rect 533682 -960 533794 480
rect 534552 354 534580 1022
rect 534878 354 534990 480
rect 534552 326 534990 354
rect 534878 -960 534990 326
rect 535380 202 535408 3060
rect 536576 2922 536604 3060
rect 536564 2916 536616 2922
rect 536564 2858 536616 2864
rect 536104 1012 536156 1018
rect 536104 954 536156 960
rect 536116 480 536144 954
rect 537680 746 537708 3060
rect 538128 1148 538180 1154
rect 538128 1090 538180 1096
rect 537208 740 537260 746
rect 537208 682 537260 688
rect 537668 740 537720 746
rect 537668 682 537720 688
rect 537220 480 537248 682
rect 535368 196 535420 202
rect 535368 138 535420 144
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538140 354 538168 1090
rect 538374 354 538486 480
rect 538140 326 538486 354
rect 538374 -960 538486 326
rect 538784 270 538812 3060
rect 539888 1358 539916 3060
rect 539876 1352 539928 1358
rect 539876 1294 539928 1300
rect 539600 672 539652 678
rect 539600 614 539652 620
rect 540900 626 540928 3060
rect 542096 678 542124 3060
rect 543214 3046 543504 3062
rect 544318 3046 544608 3074
rect 544384 876 544436 882
rect 544384 818 544436 824
rect 542084 672 542136 678
rect 539612 480 539640 614
rect 540900 598 541020 626
rect 542084 614 542136 620
rect 538772 264 538824 270
rect 538772 206 538824 212
rect 539570 -960 539682 480
rect 540428 400 540480 406
rect 540766 354 540878 480
rect 540480 348 540878 354
rect 540428 342 540878 348
rect 540440 326 540878 342
rect 540766 -960 540878 326
rect 540992 134 541020 598
rect 544396 480 544424 818
rect 541962 354 542074 480
rect 542176 468 542228 474
rect 542176 410 542228 416
rect 542188 354 542216 410
rect 541962 326 542216 354
rect 540980 128 541032 134
rect 540980 70 541032 76
rect 541962 -960 542074 326
rect 543158 82 543270 480
rect 542832 66 543270 82
rect 542820 60 543270 66
rect 542872 54 543270 60
rect 542820 2 542872 8
rect 543158 -960 543270 54
rect 544354 -960 544466 480
rect 544580 474 544608 3046
rect 545408 610 545436 3060
rect 545488 808 545540 814
rect 545488 750 545540 756
rect 545396 604 545448 610
rect 545396 546 545448 552
rect 545500 480 545528 750
rect 544568 468 544620 474
rect 544568 410 544620 416
rect 545458 -960 545570 480
rect 546420 66 546448 3060
rect 546684 3052 546736 3058
rect 546684 2994 546736 3000
rect 546696 480 546724 2994
rect 547616 882 547644 3060
rect 548734 3046 549024 3074
rect 548708 944 548760 950
rect 548708 886 548760 892
rect 547604 876 547656 882
rect 547604 818 547656 824
rect 546408 60 546460 66
rect 546408 2 546460 8
rect 546654 -960 546766 480
rect 547850 354 547962 480
rect 548720 354 548748 886
rect 548996 678 549024 3046
rect 549824 2990 549852 3060
rect 549812 2984 549864 2990
rect 549812 2926 549864 2932
rect 550928 814 550956 3060
rect 551100 1284 551152 1290
rect 551100 1226 551152 1232
rect 550916 808 550968 814
rect 550916 750 550968 756
rect 548984 672 549036 678
rect 548984 614 549036 620
rect 549046 354 549158 480
rect 547850 338 548104 354
rect 547850 332 548116 338
rect 547850 326 548064 332
rect 547850 -960 547962 326
rect 548720 326 549158 354
rect 548064 274 548116 280
rect 549046 -960 549158 326
rect 550242 354 550354 480
rect 550456 400 550508 406
rect 550242 348 550456 354
rect 550242 342 550508 348
rect 551112 354 551140 1226
rect 551438 354 551550 480
rect 550242 326 550496 342
rect 551112 326 551550 354
rect 551940 338 551968 3060
rect 553150 3058 553348 3074
rect 553150 3052 553360 3058
rect 553150 3046 553308 3052
rect 553308 2994 553360 3000
rect 553768 2916 553820 2922
rect 553768 2858 553820 2864
rect 553780 480 553808 2858
rect 550242 -960 550354 326
rect 551438 -960 551550 326
rect 551928 332 551980 338
rect 551928 274 551980 280
rect 552634 218 552746 480
rect 552634 202 552888 218
rect 552634 196 552900 202
rect 552634 190 552848 196
rect 552634 -960 552746 190
rect 552848 138 552900 144
rect 553738 -960 553850 480
rect 554240 202 554268 3060
rect 554964 740 555016 746
rect 554964 682 555016 688
rect 554976 480 555004 682
rect 554228 196 554280 202
rect 554228 138 554280 144
rect 554934 -960 555046 480
rect 555344 406 555372 3060
rect 557184 3046 557474 3074
rect 558670 3046 558868 3074
rect 562232 3120 562284 3126
rect 560484 3062 560536 3068
rect 561982 3068 562232 3074
rect 561982 3062 562284 3068
rect 556988 1352 557040 1358
rect 556988 1294 557040 1300
rect 555332 400 555384 406
rect 555332 342 555384 348
rect 556130 218 556242 480
rect 556344 264 556396 270
rect 556130 212 556344 218
rect 556130 206 556396 212
rect 556130 190 556384 206
rect 556130 -960 556242 190
rect 557000 82 557028 1294
rect 557184 270 557212 3046
rect 557172 264 557224 270
rect 557172 206 557224 212
rect 557326 82 557438 480
rect 557000 54 557438 82
rect 557326 -960 557438 54
rect 558522 82 558634 480
rect 558840 134 558868 3046
rect 559760 2922 559788 3060
rect 559748 2916 559800 2922
rect 559748 2858 559800 2864
rect 559380 536 559432 542
rect 559380 478 559432 484
rect 559392 354 559420 478
rect 559718 354 559830 480
rect 559392 326 559830 354
rect 560496 354 560524 3062
rect 561982 3046 562272 3062
rect 562980 2854 563008 3060
rect 571524 3052 571576 3058
rect 571524 2994 571576 3000
rect 568028 2984 568080 2990
rect 568028 2926 568080 2932
rect 562968 2848 563020 2854
rect 562968 2790 563020 2796
rect 565636 876 565688 882
rect 565636 818 565688 824
rect 563244 604 563296 610
rect 563244 546 563296 552
rect 563256 480 563284 546
rect 565648 480 565676 818
rect 566832 672 566884 678
rect 566832 614 566884 620
rect 566844 480 566872 614
rect 568040 480 568068 2926
rect 569132 808 569184 814
rect 569132 750 569184 756
rect 569144 480 569172 750
rect 571536 480 571564 2994
rect 575124 480 575152 3198
rect 579804 3188 579856 3194
rect 579804 3130 579856 3136
rect 578608 2916 578660 2922
rect 578608 2858 578660 2864
rect 578620 480 578648 2858
rect 579816 480 579844 3130
rect 581000 3120 581052 3126
rect 581000 3062 581052 3068
rect 581012 480 581040 3062
rect 582196 2848 582248 2854
rect 582196 2790 582248 2796
rect 582208 480 582236 2790
rect 583404 480 583432 3266
rect 560822 354 560934 480
rect 560496 326 560934 354
rect 558736 128 558788 134
rect 558522 76 558736 82
rect 558522 70 558788 76
rect 558828 128 558880 134
rect 558828 70 558880 76
rect 558522 54 558776 70
rect 558522 -960 558634 54
rect 559718 -960 559830 326
rect 560822 -960 560934 326
rect 562018 354 562130 480
rect 562232 468 562284 474
rect 562232 410 562284 416
rect 562244 354 562272 410
rect 562018 326 562272 354
rect 562018 -960 562130 326
rect 563214 -960 563326 480
rect 564410 82 564522 480
rect 564410 66 564664 82
rect 564410 60 564676 66
rect 564410 54 564624 60
rect 564410 -960 564522 54
rect 564624 2 564676 8
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 354 570410 480
rect 570298 338 570552 354
rect 570298 332 570564 338
rect 570298 326 570512 332
rect 570298 -960 570410 326
rect 570512 274 570564 280
rect 571494 -960 571606 480
rect 572690 218 572802 480
rect 573548 400 573600 406
rect 573886 354 573998 480
rect 573600 348 573998 354
rect 573548 342 573998 348
rect 573560 326 573998 342
rect 572690 202 572944 218
rect 572690 196 572956 202
rect 572690 190 572904 196
rect 572690 -960 572802 190
rect 572904 138 572956 144
rect 573886 -960 573998 326
rect 575082 -960 575194 480
rect 575940 264 575992 270
rect 576278 218 576390 480
rect 575992 212 576390 218
rect 575940 206 576390 212
rect 575952 190 576390 206
rect 576278 -960 576390 190
rect 577136 128 577188 134
rect 577382 82 577494 480
rect 577188 76 577494 82
rect 577136 70 577494 76
rect 577148 54 577494 70
rect 577382 -960 577494 54
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 2778 697312 2834 697368
rect 581642 697176 581698 697232
rect 581642 691464 581698 691520
rect 2778 690784 2834 690840
rect 2778 684256 2834 684312
rect 582378 683848 582434 683904
rect 582378 678408 582434 678464
rect 2778 678000 2834 678056
rect 2778 671200 2834 671256
rect 582378 670656 582434 670712
rect 582378 665352 582434 665408
rect 2778 665216 2834 665272
rect 2778 658144 2834 658200
rect 582378 657328 582434 657384
rect 2778 652432 2834 652488
rect 582378 652296 582434 652352
rect 2778 645088 2834 645144
rect 581642 644000 581698 644056
rect 2778 639648 2834 639704
rect 581642 639240 581698 639296
rect 2778 632032 2834 632088
rect 582378 630808 582434 630864
rect 2778 626864 2834 626920
rect 582378 626184 582434 626240
rect 2778 619112 2834 619168
rect 581642 617480 581698 617536
rect 2778 613944 2834 614000
rect 581642 613128 581698 613184
rect 2778 606056 2834 606112
rect 581642 604152 581698 604208
rect 2778 601296 2834 601352
rect 581642 600072 581698 600128
rect 1582 593000 1638 593056
rect 581642 590960 581698 591016
rect 1582 588512 1638 588568
rect 581642 587016 581698 587072
rect 2042 579944 2098 580000
rect 581642 577632 581698 577688
rect 2042 575728 2098 575784
rect 581642 573960 581698 574016
rect 1490 566888 1546 566944
rect 582378 564304 582434 564360
rect 1490 562944 1546 563000
rect 582378 560904 582434 560960
rect 1490 553832 1546 553888
rect 581642 551112 581698 551168
rect 1490 550160 1546 550216
rect 581642 547712 581698 547768
rect 1398 540776 1454 540832
rect 582378 537784 582434 537840
rect 1398 537376 1454 537432
rect 582378 534792 582434 534848
rect 1490 527856 1546 527912
rect 1490 524592 1546 524648
rect 582378 524456 582434 524512
rect 582378 521736 582434 521792
rect 1582 514800 1638 514856
rect 1582 511808 1638 511864
rect 582378 511264 582434 511320
rect 582378 508680 582434 508736
rect 1582 501744 1638 501800
rect 1582 499024 1638 499080
rect 581642 497936 581698 497992
rect 581642 495624 581698 495680
rect 1582 488688 1638 488744
rect 1582 486240 1638 486296
rect 582378 484608 582434 484664
rect 582378 482568 582434 482624
rect 2778 475632 2834 475688
rect 2778 473456 2834 473512
rect 581642 471416 581698 471472
rect 581642 469512 581698 469568
rect 1582 462576 1638 462632
rect 1582 460672 1638 460728
rect 581642 458088 581698 458144
rect 581642 456456 581698 456512
rect 2778 449520 2834 449576
rect 2778 447888 2834 447944
rect 2778 436600 2834 436656
rect 2778 435104 2834 435160
rect 2778 423544 2834 423600
rect 2778 422320 2834 422376
rect 1306 294344 1362 294400
rect 1306 293120 1362 293176
rect 2778 281560 2834 281616
rect 2778 280064 2834 280120
rect 1306 268776 1362 268832
rect 1306 267144 1362 267200
rect 582378 260480 582434 260536
rect 582378 258848 582434 258904
rect 1306 255992 1362 256048
rect 1306 254088 1362 254144
rect 580906 247016 580962 247072
rect 580906 245520 580962 245576
rect 2778 243208 2834 243264
rect 2778 241032 2834 241088
rect 582378 234368 582434 234424
rect 582378 232328 582434 232384
rect 2778 230560 2834 230616
rect 2778 227976 2834 228032
rect 580906 220904 580962 220960
rect 580906 219000 580962 219056
rect 2778 217640 2834 217696
rect 2778 214920 2834 214976
rect 582378 208256 582434 208312
rect 582378 205672 582434 205728
rect 2778 204856 2834 204912
rect 2778 201864 2834 201920
rect 580906 194656 580962 194712
rect 580906 192480 580962 192536
rect 1306 192072 1362 192128
rect 1306 188808 1362 188864
rect 580906 182416 580962 182472
rect 2778 179288 2834 179344
rect 580906 179152 580962 179208
rect 2778 175888 2834 175944
rect 580906 168544 580962 168600
rect 2778 166504 2834 166560
rect 580906 165824 580962 165880
rect 2778 162832 2834 162888
rect 580906 156304 580962 156360
rect 1306 153720 1362 153776
rect 580906 152632 580962 152688
rect 1306 149776 1362 149832
rect 580906 142568 580962 142624
rect 570 140936 626 140992
rect 580906 139304 580962 139360
rect 570 136720 626 136776
rect 580906 130192 580962 130248
rect 754 128152 810 128208
rect 580906 125976 580962 126032
rect 754 123664 810 123720
rect 579894 116320 579950 116376
rect 1306 115368 1362 115424
rect 579894 112784 579950 112840
rect 1306 110608 1362 110664
rect 580906 103536 580962 103592
rect 1582 102584 1638 102640
rect 580906 99456 580962 99512
rect 1582 97552 1638 97608
rect 580906 90208 580962 90264
rect 1582 89800 1638 89856
rect 580906 86128 580962 86184
rect 1582 84632 1638 84688
rect 579894 77288 579950 77344
rect 1582 77016 1638 77072
rect 579894 72936 579950 72992
rect 1582 71576 1638 71632
rect 1490 64232 1546 64288
rect 580906 64096 580962 64152
rect 580906 59608 580962 59664
rect 1490 58520 1546 58576
rect 2042 51448 2098 51504
rect 580906 51040 580962 51096
rect 580906 46280 580962 46336
rect 2042 45464 2098 45520
rect 2042 38664 2098 38720
rect 580906 37984 580962 38040
rect 580906 33088 580962 33144
rect 2042 32408 2098 32464
rect 1490 25880 1546 25936
rect 580906 24928 580962 24984
rect 580906 19760 580962 19816
rect 1490 19352 1546 19408
rect 2042 13096 2098 13152
rect 579894 12688 579950 12744
rect 579894 6568 579950 6624
rect 2042 6432 2098 6488
rect 70214 3884 70216 3904
rect 70216 3884 70268 3904
rect 70268 3884 70270 3904
rect 70214 3848 70270 3884
rect 73618 3848 73674 3904
rect 5446 312 5502 368
rect 6274 40 6330 96
rect 12162 448 12218 504
rect 13726 176 13782 232
rect 23938 312 23994 368
rect 25042 40 25098 96
rect 25686 312 25742 368
rect 28906 584 28962 640
rect 30838 448 30894 504
rect 31942 176 31998 232
rect 37002 176 37058 232
rect 42706 312 42762 368
rect 46294 584 46350 640
rect 46846 40 46902 96
rect 54022 176 54078 232
rect 62854 40 62910 96
<< metal3 >>
rect -960 697370 480 697460
rect 2773 697370 2839 697373
rect -960 697368 2839 697370
rect -960 697312 2778 697368
rect 2834 697312 2839 697368
rect -960 697310 2839 697312
rect -960 697220 480 697310
rect 2773 697307 2839 697310
rect 581637 697234 581703 697237
rect 583520 697234 584960 697324
rect 581637 697232 584960 697234
rect 581637 697176 581642 697232
rect 581698 697176 584960 697232
rect 581637 697174 584960 697176
rect 581637 697171 581703 697174
rect 583520 697084 584960 697174
rect 581637 691522 581703 691525
rect 580796 691520 581703 691522
rect 580796 691464 581642 691520
rect 581698 691464 581703 691520
rect 580796 691462 581703 691464
rect 581637 691459 581703 691462
rect 2773 690842 2839 690845
rect 2773 690840 3220 690842
rect 2773 690784 2778 690840
rect 2834 690784 3220 690840
rect 2773 690782 3220 690784
rect 2773 690779 2839 690782
rect -960 684314 480 684404
rect 2773 684314 2839 684317
rect -960 684312 2839 684314
rect -960 684256 2778 684312
rect 2834 684256 2839 684312
rect -960 684254 2839 684256
rect -960 684164 480 684254
rect 2773 684251 2839 684254
rect 582373 683906 582439 683909
rect 583520 683906 584960 683996
rect 582373 683904 584960 683906
rect 582373 683848 582378 683904
rect 582434 683848 584960 683904
rect 582373 683846 584960 683848
rect 582373 683843 582439 683846
rect 583520 683756 584960 683846
rect 582373 678466 582439 678469
rect 580796 678464 582439 678466
rect 580796 678408 582378 678464
rect 582434 678408 582439 678464
rect 580796 678406 582439 678408
rect 582373 678403 582439 678406
rect 2773 678058 2839 678061
rect 2773 678056 3220 678058
rect 2773 678000 2778 678056
rect 2834 678000 3220 678056
rect 2773 677998 3220 678000
rect 2773 677995 2839 677998
rect -960 671258 480 671348
rect 2773 671258 2839 671261
rect -960 671256 2839 671258
rect -960 671200 2778 671256
rect 2834 671200 2839 671256
rect -960 671198 2839 671200
rect -960 671108 480 671198
rect 2773 671195 2839 671198
rect 582373 670714 582439 670717
rect 583520 670714 584960 670804
rect 582373 670712 584960 670714
rect 582373 670656 582378 670712
rect 582434 670656 584960 670712
rect 582373 670654 584960 670656
rect 582373 670651 582439 670654
rect 583520 670564 584960 670654
rect 582373 665410 582439 665413
rect 580796 665408 582439 665410
rect 580796 665352 582378 665408
rect 582434 665352 582439 665408
rect 580796 665350 582439 665352
rect 582373 665347 582439 665350
rect 2773 665274 2839 665277
rect 2773 665272 3220 665274
rect 2773 665216 2778 665272
rect 2834 665216 3220 665272
rect 2773 665214 3220 665216
rect 2773 665211 2839 665214
rect -960 658202 480 658292
rect 2773 658202 2839 658205
rect -960 658200 2839 658202
rect -960 658144 2778 658200
rect 2834 658144 2839 658200
rect -960 658142 2839 658144
rect -960 658052 480 658142
rect 2773 658139 2839 658142
rect 582373 657386 582439 657389
rect 583520 657386 584960 657476
rect 582373 657384 584960 657386
rect 582373 657328 582378 657384
rect 582434 657328 584960 657384
rect 582373 657326 584960 657328
rect 582373 657323 582439 657326
rect 583520 657236 584960 657326
rect 2773 652490 2839 652493
rect 2773 652488 3220 652490
rect 2773 652432 2778 652488
rect 2834 652432 3220 652488
rect 2773 652430 3220 652432
rect 2773 652427 2839 652430
rect 582373 652354 582439 652357
rect 580796 652352 582439 652354
rect 580796 652296 582378 652352
rect 582434 652296 582439 652352
rect 580796 652294 582439 652296
rect 582373 652291 582439 652294
rect -960 645146 480 645236
rect 2773 645146 2839 645149
rect -960 645144 2839 645146
rect -960 645088 2778 645144
rect 2834 645088 2839 645144
rect -960 645086 2839 645088
rect -960 644996 480 645086
rect 2773 645083 2839 645086
rect 581637 644058 581703 644061
rect 583520 644058 584960 644148
rect 581637 644056 584960 644058
rect 581637 644000 581642 644056
rect 581698 644000 584960 644056
rect 581637 643998 584960 644000
rect 581637 643995 581703 643998
rect 583520 643908 584960 643998
rect 2773 639706 2839 639709
rect 2773 639704 3220 639706
rect 2773 639648 2778 639704
rect 2834 639648 3220 639704
rect 2773 639646 3220 639648
rect 2773 639643 2839 639646
rect 581637 639298 581703 639301
rect 580796 639296 581703 639298
rect 580796 639240 581642 639296
rect 581698 639240 581703 639296
rect 580796 639238 581703 639240
rect 581637 639235 581703 639238
rect -960 632090 480 632180
rect 2773 632090 2839 632093
rect -960 632088 2839 632090
rect -960 632032 2778 632088
rect 2834 632032 2839 632088
rect -960 632030 2839 632032
rect -960 631940 480 632030
rect 2773 632027 2839 632030
rect 582373 630866 582439 630869
rect 583520 630866 584960 630956
rect 582373 630864 584960 630866
rect 582373 630808 582378 630864
rect 582434 630808 584960 630864
rect 582373 630806 584960 630808
rect 582373 630803 582439 630806
rect 583520 630716 584960 630806
rect 2773 626922 2839 626925
rect 2773 626920 3220 626922
rect 2773 626864 2778 626920
rect 2834 626864 3220 626920
rect 2773 626862 3220 626864
rect 2773 626859 2839 626862
rect 582373 626242 582439 626245
rect 580796 626240 582439 626242
rect 580796 626184 582378 626240
rect 582434 626184 582439 626240
rect 580796 626182 582439 626184
rect 582373 626179 582439 626182
rect -960 619170 480 619260
rect 2773 619170 2839 619173
rect -960 619168 2839 619170
rect -960 619112 2778 619168
rect 2834 619112 2839 619168
rect -960 619110 2839 619112
rect -960 619020 480 619110
rect 2773 619107 2839 619110
rect 581637 617538 581703 617541
rect 583520 617538 584960 617628
rect 581637 617536 584960 617538
rect 581637 617480 581642 617536
rect 581698 617480 584960 617536
rect 581637 617478 584960 617480
rect 581637 617475 581703 617478
rect 583520 617388 584960 617478
rect 2773 614002 2839 614005
rect 2773 614000 3220 614002
rect 2773 613944 2778 614000
rect 2834 613944 3220 614000
rect 2773 613942 3220 613944
rect 2773 613939 2839 613942
rect 581637 613186 581703 613189
rect 580796 613184 581703 613186
rect 580796 613128 581642 613184
rect 581698 613128 581703 613184
rect 580796 613126 581703 613128
rect 581637 613123 581703 613126
rect -960 606114 480 606204
rect 2773 606114 2839 606117
rect -960 606112 2839 606114
rect -960 606056 2778 606112
rect 2834 606056 2839 606112
rect -960 606054 2839 606056
rect -960 605964 480 606054
rect 2773 606051 2839 606054
rect 581637 604210 581703 604213
rect 583520 604210 584960 604300
rect 581637 604208 584960 604210
rect 581637 604152 581642 604208
rect 581698 604152 584960 604208
rect 581637 604150 584960 604152
rect 581637 604147 581703 604150
rect 583520 604060 584960 604150
rect 2773 601354 2839 601357
rect 2773 601352 3220 601354
rect 2773 601296 2778 601352
rect 2834 601296 3220 601352
rect 2773 601294 3220 601296
rect 2773 601291 2839 601294
rect 581637 600130 581703 600133
rect 580796 600128 581703 600130
rect 580796 600072 581642 600128
rect 581698 600072 581703 600128
rect 580796 600070 581703 600072
rect 581637 600067 581703 600070
rect -960 593058 480 593148
rect 1577 593058 1643 593061
rect -960 593056 1643 593058
rect -960 593000 1582 593056
rect 1638 593000 1643 593056
rect -960 592998 1643 593000
rect -960 592908 480 592998
rect 1577 592995 1643 592998
rect 581637 591018 581703 591021
rect 583520 591018 584960 591108
rect 581637 591016 584960 591018
rect 581637 590960 581642 591016
rect 581698 590960 584960 591016
rect 581637 590958 584960 590960
rect 581637 590955 581703 590958
rect 583520 590868 584960 590958
rect 1577 588570 1643 588573
rect 1577 588568 3220 588570
rect 1577 588512 1582 588568
rect 1638 588512 3220 588568
rect 1577 588510 3220 588512
rect 1577 588507 1643 588510
rect 581637 587074 581703 587077
rect 580796 587072 581703 587074
rect 580796 587016 581642 587072
rect 581698 587016 581703 587072
rect 580796 587014 581703 587016
rect 581637 587011 581703 587014
rect -960 580002 480 580092
rect 2037 580002 2103 580005
rect -960 580000 2103 580002
rect -960 579944 2042 580000
rect 2098 579944 2103 580000
rect -960 579942 2103 579944
rect -960 579852 480 579942
rect 2037 579939 2103 579942
rect 581637 577690 581703 577693
rect 583520 577690 584960 577780
rect 581637 577688 584960 577690
rect 581637 577632 581642 577688
rect 581698 577632 584960 577688
rect 581637 577630 584960 577632
rect 581637 577627 581703 577630
rect 583520 577540 584960 577630
rect 2037 575786 2103 575789
rect 2037 575784 3220 575786
rect 2037 575728 2042 575784
rect 2098 575728 3220 575784
rect 2037 575726 3220 575728
rect 2037 575723 2103 575726
rect 581637 574018 581703 574021
rect 580796 574016 581703 574018
rect 580796 573960 581642 574016
rect 581698 573960 581703 574016
rect 580796 573958 581703 573960
rect 581637 573955 581703 573958
rect -960 566946 480 567036
rect 1485 566946 1551 566949
rect -960 566944 1551 566946
rect -960 566888 1490 566944
rect 1546 566888 1551 566944
rect -960 566886 1551 566888
rect -960 566796 480 566886
rect 1485 566883 1551 566886
rect 582373 564362 582439 564365
rect 583520 564362 584960 564452
rect 582373 564360 584960 564362
rect 582373 564304 582378 564360
rect 582434 564304 584960 564360
rect 582373 564302 584960 564304
rect 582373 564299 582439 564302
rect 583520 564212 584960 564302
rect 1485 563002 1551 563005
rect 1485 563000 3220 563002
rect 1485 562944 1490 563000
rect 1546 562944 3220 563000
rect 1485 562942 3220 562944
rect 1485 562939 1551 562942
rect 582373 560962 582439 560965
rect 580796 560960 582439 560962
rect 580796 560904 582378 560960
rect 582434 560904 582439 560960
rect 580796 560902 582439 560904
rect 582373 560899 582439 560902
rect -960 553890 480 553980
rect 1485 553890 1551 553893
rect -960 553888 1551 553890
rect -960 553832 1490 553888
rect 1546 553832 1551 553888
rect -960 553830 1551 553832
rect -960 553740 480 553830
rect 1485 553827 1551 553830
rect 581637 551170 581703 551173
rect 583520 551170 584960 551260
rect 581637 551168 584960 551170
rect 581637 551112 581642 551168
rect 581698 551112 584960 551168
rect 581637 551110 584960 551112
rect 581637 551107 581703 551110
rect 583520 551020 584960 551110
rect 1485 550218 1551 550221
rect 1485 550216 3220 550218
rect 1485 550160 1490 550216
rect 1546 550160 3220 550216
rect 1485 550158 3220 550160
rect 1485 550155 1551 550158
rect 581637 547770 581703 547773
rect 580796 547768 581703 547770
rect 580796 547712 581642 547768
rect 581698 547712 581703 547768
rect 580796 547710 581703 547712
rect 581637 547707 581703 547710
rect -960 540834 480 540924
rect 1393 540834 1459 540837
rect -960 540832 1459 540834
rect -960 540776 1398 540832
rect 1454 540776 1459 540832
rect -960 540774 1459 540776
rect -960 540684 480 540774
rect 1393 540771 1459 540774
rect 582373 537842 582439 537845
rect 583520 537842 584960 537932
rect 582373 537840 584960 537842
rect 582373 537784 582378 537840
rect 582434 537784 584960 537840
rect 582373 537782 584960 537784
rect 582373 537779 582439 537782
rect 583520 537692 584960 537782
rect 1393 537434 1459 537437
rect 1393 537432 3220 537434
rect 1393 537376 1398 537432
rect 1454 537376 3220 537432
rect 1393 537374 3220 537376
rect 1393 537371 1459 537374
rect 582373 534850 582439 534853
rect 580796 534848 582439 534850
rect 580796 534792 582378 534848
rect 582434 534792 582439 534848
rect 580796 534790 582439 534792
rect 582373 534787 582439 534790
rect -960 527914 480 528004
rect 1485 527914 1551 527917
rect -960 527912 1551 527914
rect -960 527856 1490 527912
rect 1546 527856 1551 527912
rect -960 527854 1551 527856
rect -960 527764 480 527854
rect 1485 527851 1551 527854
rect 1485 524650 1551 524653
rect 1485 524648 3220 524650
rect 1485 524592 1490 524648
rect 1546 524592 3220 524648
rect 1485 524590 3220 524592
rect 1485 524587 1551 524590
rect 582373 524514 582439 524517
rect 583520 524514 584960 524604
rect 582373 524512 584960 524514
rect 582373 524456 582378 524512
rect 582434 524456 584960 524512
rect 582373 524454 584960 524456
rect 582373 524451 582439 524454
rect 583520 524364 584960 524454
rect 582373 521794 582439 521797
rect 580796 521792 582439 521794
rect 580796 521736 582378 521792
rect 582434 521736 582439 521792
rect 580796 521734 582439 521736
rect 582373 521731 582439 521734
rect -960 514858 480 514948
rect 1577 514858 1643 514861
rect -960 514856 1643 514858
rect -960 514800 1582 514856
rect 1638 514800 1643 514856
rect -960 514798 1643 514800
rect -960 514708 480 514798
rect 1577 514795 1643 514798
rect 1577 511866 1643 511869
rect 1577 511864 3220 511866
rect 1577 511808 1582 511864
rect 1638 511808 3220 511864
rect 1577 511806 3220 511808
rect 1577 511803 1643 511806
rect 582373 511322 582439 511325
rect 583520 511322 584960 511412
rect 582373 511320 584960 511322
rect 582373 511264 582378 511320
rect 582434 511264 584960 511320
rect 582373 511262 584960 511264
rect 582373 511259 582439 511262
rect 583520 511172 584960 511262
rect 582373 508738 582439 508741
rect 580796 508736 582439 508738
rect 580796 508680 582378 508736
rect 582434 508680 582439 508736
rect 580796 508678 582439 508680
rect 582373 508675 582439 508678
rect -960 501802 480 501892
rect 1577 501802 1643 501805
rect -960 501800 1643 501802
rect -960 501744 1582 501800
rect 1638 501744 1643 501800
rect -960 501742 1643 501744
rect -960 501652 480 501742
rect 1577 501739 1643 501742
rect 1577 499082 1643 499085
rect 1577 499080 3220 499082
rect 1577 499024 1582 499080
rect 1638 499024 3220 499080
rect 1577 499022 3220 499024
rect 1577 499019 1643 499022
rect 581637 497994 581703 497997
rect 583520 497994 584960 498084
rect 581637 497992 584960 497994
rect 581637 497936 581642 497992
rect 581698 497936 584960 497992
rect 581637 497934 584960 497936
rect 581637 497931 581703 497934
rect 583520 497844 584960 497934
rect 581637 495682 581703 495685
rect 580796 495680 581703 495682
rect 580796 495624 581642 495680
rect 581698 495624 581703 495680
rect 580796 495622 581703 495624
rect 581637 495619 581703 495622
rect -960 488746 480 488836
rect 1577 488746 1643 488749
rect -960 488744 1643 488746
rect -960 488688 1582 488744
rect 1638 488688 1643 488744
rect -960 488686 1643 488688
rect -960 488596 480 488686
rect 1577 488683 1643 488686
rect 1577 486298 1643 486301
rect 1577 486296 3220 486298
rect 1577 486240 1582 486296
rect 1638 486240 3220 486296
rect 1577 486238 3220 486240
rect 1577 486235 1643 486238
rect 582373 484666 582439 484669
rect 583520 484666 584960 484756
rect 582373 484664 584960 484666
rect 582373 484608 582378 484664
rect 582434 484608 584960 484664
rect 582373 484606 584960 484608
rect 582373 484603 582439 484606
rect 583520 484516 584960 484606
rect 582373 482626 582439 482629
rect 580796 482624 582439 482626
rect 580796 482568 582378 482624
rect 582434 482568 582439 482624
rect 580796 482566 582439 482568
rect 582373 482563 582439 482566
rect -960 475690 480 475780
rect 2773 475690 2839 475693
rect -960 475688 2839 475690
rect -960 475632 2778 475688
rect 2834 475632 2839 475688
rect -960 475630 2839 475632
rect -960 475540 480 475630
rect 2773 475627 2839 475630
rect 2773 473514 2839 473517
rect 2773 473512 3220 473514
rect 2773 473456 2778 473512
rect 2834 473456 3220 473512
rect 2773 473454 3220 473456
rect 2773 473451 2839 473454
rect 581637 471474 581703 471477
rect 583520 471474 584960 471564
rect 581637 471472 584960 471474
rect 581637 471416 581642 471472
rect 581698 471416 584960 471472
rect 581637 471414 584960 471416
rect 581637 471411 581703 471414
rect 583520 471324 584960 471414
rect 581637 469570 581703 469573
rect 580796 469568 581703 469570
rect 580796 469512 581642 469568
rect 581698 469512 581703 469568
rect 580796 469510 581703 469512
rect 581637 469507 581703 469510
rect -960 462634 480 462724
rect 1577 462634 1643 462637
rect -960 462632 1643 462634
rect -960 462576 1582 462632
rect 1638 462576 1643 462632
rect -960 462574 1643 462576
rect -960 462484 480 462574
rect 1577 462571 1643 462574
rect 1577 460730 1643 460733
rect 1577 460728 3220 460730
rect 1577 460672 1582 460728
rect 1638 460672 3220 460728
rect 1577 460670 3220 460672
rect 1577 460667 1643 460670
rect 581637 458146 581703 458149
rect 583520 458146 584960 458236
rect 581637 458144 584960 458146
rect 581637 458088 581642 458144
rect 581698 458088 584960 458144
rect 581637 458086 584960 458088
rect 581637 458083 581703 458086
rect 583520 457996 584960 458086
rect 581637 456514 581703 456517
rect 580796 456512 581703 456514
rect 580796 456456 581642 456512
rect 581698 456456 581703 456512
rect 580796 456454 581703 456456
rect 581637 456451 581703 456454
rect -960 449578 480 449668
rect 2773 449578 2839 449581
rect -960 449576 2839 449578
rect -960 449520 2778 449576
rect 2834 449520 2839 449576
rect -960 449518 2839 449520
rect -960 449428 480 449518
rect 2773 449515 2839 449518
rect 2773 447946 2839 447949
rect 2773 447944 3220 447946
rect 2773 447888 2778 447944
rect 2834 447888 3220 447944
rect 2773 447886 3220 447888
rect 2773 447883 2839 447886
rect 583520 444818 584960 444908
rect 583342 444758 584960 444818
rect 583342 444682 583402 444758
rect 583520 444682 584960 444758
rect 583342 444668 584960 444682
rect 583342 444622 583586 444668
rect 583526 444138 583586 444622
rect 580766 444078 583586 444138
rect 580766 443428 580826 444078
rect -960 436658 480 436748
rect 2773 436658 2839 436661
rect -960 436656 2839 436658
rect -960 436600 2778 436656
rect 2834 436600 2839 436656
rect -960 436598 2839 436600
rect -960 436508 480 436598
rect 2773 436595 2839 436598
rect 2773 435162 2839 435165
rect 2773 435160 3220 435162
rect 2773 435104 2778 435160
rect 2834 435104 3220 435160
rect 2773 435102 3220 435104
rect 2773 435099 2839 435102
rect 583520 431626 584960 431716
rect 583342 431566 584960 431626
rect 583342 431490 583402 431566
rect 583520 431490 584960 431566
rect 583342 431476 584960 431490
rect 583342 431430 583586 431476
rect 583526 431082 583586 431430
rect 580766 431022 583586 431082
rect 580766 430372 580826 431022
rect -960 423602 480 423692
rect 2773 423602 2839 423605
rect -960 423600 2839 423602
rect -960 423544 2778 423600
rect 2834 423544 2839 423600
rect -960 423542 2839 423544
rect -960 423452 480 423542
rect 2773 423539 2839 423542
rect 2773 422378 2839 422381
rect 2773 422376 3220 422378
rect 2773 422320 2778 422376
rect 2834 422320 3220 422376
rect 2773 422318 3220 422320
rect 2773 422315 2839 422318
rect 583520 418298 584960 418388
rect 583342 418238 584960 418298
rect 583342 418162 583402 418238
rect 583520 418162 584960 418238
rect 583342 418148 584960 418162
rect 583342 418102 583586 418148
rect 583526 417754 583586 418102
rect 580766 417694 583586 417754
rect 580766 417316 580826 417694
rect -960 410546 480 410636
rect -960 410486 3250 410546
rect -960 410396 480 410486
rect 3190 409564 3250 410486
rect 583520 404970 584960 405060
rect 580766 404910 584960 404970
rect 580766 404260 580826 404910
rect 583520 404820 584960 404910
rect -960 397490 480 397580
rect -960 397430 3250 397490
rect -960 397340 480 397430
rect 3190 396780 3250 397430
rect 583520 391778 584960 391868
rect 580766 391718 584960 391778
rect 580766 391204 580826 391718
rect 583520 391628 584960 391718
rect -960 384434 480 384524
rect -960 384374 3250 384434
rect -960 384284 480 384374
rect 3190 383996 3250 384374
rect 583520 378450 584960 378540
rect 580766 378390 584960 378450
rect 580766 378148 580826 378390
rect 583520 378300 584960 378390
rect -960 371378 480 371468
rect -960 371318 3250 371378
rect -960 371228 480 371318
rect 3190 371212 3250 371318
rect 583520 365122 584960 365212
rect 580796 365062 584960 365122
rect 583520 364972 584960 365062
rect -960 358458 480 358548
rect -960 358398 3220 358458
rect -960 358308 480 358398
rect 583520 351930 584960 352020
rect 580796 351870 584960 351930
rect 583520 351780 584960 351870
rect -960 345402 480 345492
rect 1534 345478 3220 345538
rect 1534 345402 1594 345478
rect -960 345342 1594 345402
rect -960 345252 480 345342
rect 580766 338602 580826 338844
rect 583520 338602 584960 338692
rect 580766 338542 584960 338602
rect 583520 338452 584960 338542
rect -960 332346 480 332436
rect 3190 332346 3250 332724
rect -960 332286 3250 332346
rect -960 332196 480 332286
rect 580766 325274 580826 325788
rect 583520 325274 584960 325364
rect 580766 325214 584960 325274
rect 583520 325124 584960 325214
rect -960 319290 480 319380
rect 3190 319290 3250 319940
rect -960 319230 3250 319290
rect -960 319140 480 319230
rect 580766 312082 580826 312732
rect 583520 312082 584960 312172
rect 580766 312022 584960 312082
rect 583520 311932 584960 312022
rect -960 306234 480 306324
rect 3190 306234 3250 307156
rect -960 306174 3250 306234
rect -960 306084 480 306174
rect 580766 299298 580826 299676
rect 580766 299238 583586 299298
rect 583526 298890 583586 299238
rect 583342 298844 583586 298890
rect 583342 298830 584960 298844
rect 583342 298754 583402 298830
rect 583520 298754 584960 298830
rect 583342 298694 584960 298754
rect 583520 298604 584960 298694
rect 1301 294402 1367 294405
rect 1301 294400 3220 294402
rect 1301 294344 1306 294400
rect 1362 294344 3220 294400
rect 1301 294342 3220 294344
rect 1301 294339 1367 294342
rect -960 293178 480 293268
rect 1301 293178 1367 293181
rect -960 293176 1367 293178
rect -960 293120 1306 293176
rect 1362 293120 1367 293176
rect -960 293118 1367 293120
rect -960 293028 480 293118
rect 1301 293115 1367 293118
rect 580766 285970 580826 286620
rect 580766 285910 583586 285970
rect 583526 285562 583586 285910
rect 583342 285516 583586 285562
rect 583342 285502 584960 285516
rect 583342 285426 583402 285502
rect 583520 285426 584960 285502
rect 583342 285366 584960 285426
rect 583520 285276 584960 285366
rect 2773 281618 2839 281621
rect 2773 281616 3220 281618
rect 2773 281560 2778 281616
rect 2834 281560 3220 281616
rect 2773 281558 3220 281560
rect 2773 281555 2839 281558
rect -960 280122 480 280212
rect 2773 280122 2839 280125
rect -960 280120 2839 280122
rect -960 280064 2778 280120
rect 2834 280064 2839 280120
rect -960 280062 2839 280064
rect -960 279972 480 280062
rect 2773 280059 2839 280062
rect 580766 272914 580826 273564
rect 580766 272854 583586 272914
rect 583526 272370 583586 272854
rect 583342 272324 583586 272370
rect 583342 272310 584960 272324
rect 583342 272234 583402 272310
rect 583520 272234 584960 272310
rect 583342 272174 584960 272234
rect 583520 272084 584960 272174
rect 1301 268834 1367 268837
rect 1301 268832 3220 268834
rect 1301 268776 1306 268832
rect 1362 268776 3220 268832
rect 1301 268774 3220 268776
rect 1301 268771 1367 268774
rect -960 267202 480 267292
rect 1301 267202 1367 267205
rect -960 267200 1367 267202
rect -960 267144 1306 267200
rect 1362 267144 1367 267200
rect -960 267142 1367 267144
rect -960 267052 480 267142
rect 1301 267139 1367 267142
rect 582373 260538 582439 260541
rect 580796 260536 582439 260538
rect 580796 260480 582378 260536
rect 582434 260480 582439 260536
rect 580796 260478 582439 260480
rect 582373 260475 582439 260478
rect 582373 258906 582439 258909
rect 583520 258906 584960 258996
rect 582373 258904 584960 258906
rect 582373 258848 582378 258904
rect 582434 258848 584960 258904
rect 582373 258846 584960 258848
rect 582373 258843 582439 258846
rect 583520 258756 584960 258846
rect 1301 256050 1367 256053
rect 1301 256048 3220 256050
rect 1301 255992 1306 256048
rect 1362 255992 3220 256048
rect 1301 255990 3220 255992
rect 1301 255987 1367 255990
rect -960 254146 480 254236
rect 1301 254146 1367 254149
rect -960 254144 1367 254146
rect -960 254088 1306 254144
rect 1362 254088 1367 254144
rect -960 254086 1367 254088
rect -960 253996 480 254086
rect 1301 254083 1367 254086
rect 580766 247074 580826 247452
rect 580901 247074 580967 247077
rect 580766 247072 580967 247074
rect 580766 247016 580906 247072
rect 580962 247016 580967 247072
rect 580766 247014 580967 247016
rect 580901 247011 580967 247014
rect 580901 245578 580967 245581
rect 583520 245578 584960 245668
rect 580901 245576 584960 245578
rect 580901 245520 580906 245576
rect 580962 245520 584960 245576
rect 580901 245518 584960 245520
rect 580901 245515 580967 245518
rect 583520 245428 584960 245518
rect 2773 243266 2839 243269
rect 2773 243264 3220 243266
rect 2773 243208 2778 243264
rect 2834 243208 3220 243264
rect 2773 243206 3220 243208
rect 2773 243203 2839 243206
rect -960 241090 480 241180
rect 2773 241090 2839 241093
rect -960 241088 2839 241090
rect -960 241032 2778 241088
rect 2834 241032 2839 241088
rect -960 241030 2839 241032
rect -960 240940 480 241030
rect 2773 241027 2839 241030
rect 582373 234426 582439 234429
rect 580796 234424 582439 234426
rect 580796 234368 582378 234424
rect 582434 234368 582439 234424
rect 580796 234366 582439 234368
rect 582373 234363 582439 234366
rect 582373 232386 582439 232389
rect 583520 232386 584960 232476
rect 582373 232384 584960 232386
rect 582373 232328 582378 232384
rect 582434 232328 584960 232384
rect 582373 232326 584960 232328
rect 582373 232323 582439 232326
rect 583520 232236 584960 232326
rect 2773 230618 2839 230621
rect 2773 230616 3220 230618
rect 2773 230560 2778 230616
rect 2834 230560 3220 230616
rect 2773 230558 3220 230560
rect 2773 230555 2839 230558
rect -960 228034 480 228124
rect 2773 228034 2839 228037
rect -960 228032 2839 228034
rect -960 227976 2778 228032
rect 2834 227976 2839 228032
rect -960 227974 2839 227976
rect -960 227884 480 227974
rect 2773 227971 2839 227974
rect 580766 220962 580826 221340
rect 580901 220962 580967 220965
rect 580766 220960 580967 220962
rect 580766 220904 580906 220960
rect 580962 220904 580967 220960
rect 580766 220902 580967 220904
rect 580901 220899 580967 220902
rect 580901 219058 580967 219061
rect 583520 219058 584960 219148
rect 580901 219056 584960 219058
rect 580901 219000 580906 219056
rect 580962 219000 584960 219056
rect 580901 218998 584960 219000
rect 580901 218995 580967 218998
rect 583520 218908 584960 218998
rect 2773 217698 2839 217701
rect 2773 217696 3220 217698
rect 2773 217640 2778 217696
rect 2834 217640 3220 217696
rect 2773 217638 3220 217640
rect 2773 217635 2839 217638
rect -960 214978 480 215068
rect 2773 214978 2839 214981
rect -960 214976 2839 214978
rect -960 214920 2778 214976
rect 2834 214920 2839 214976
rect -960 214918 2839 214920
rect -960 214828 480 214918
rect 2773 214915 2839 214918
rect 582373 208314 582439 208317
rect 580796 208312 582439 208314
rect 580796 208256 582378 208312
rect 582434 208256 582439 208312
rect 580796 208254 582439 208256
rect 582373 208251 582439 208254
rect 582373 205730 582439 205733
rect 583520 205730 584960 205820
rect 582373 205728 584960 205730
rect 582373 205672 582378 205728
rect 582434 205672 584960 205728
rect 582373 205670 584960 205672
rect 582373 205667 582439 205670
rect 583520 205580 584960 205670
rect 2773 204914 2839 204917
rect 2773 204912 3220 204914
rect 2773 204856 2778 204912
rect 2834 204856 3220 204912
rect 2773 204854 3220 204856
rect 2773 204851 2839 204854
rect -960 201922 480 202012
rect 2773 201922 2839 201925
rect -960 201920 2839 201922
rect -960 201864 2778 201920
rect 2834 201864 2839 201920
rect -960 201862 2839 201864
rect -960 201772 480 201862
rect 2773 201859 2839 201862
rect 580766 194714 580826 195228
rect 580901 194714 580967 194717
rect 580766 194712 580967 194714
rect 580766 194656 580906 194712
rect 580962 194656 580967 194712
rect 580766 194654 580967 194656
rect 580901 194651 580967 194654
rect 580901 192538 580967 192541
rect 583520 192538 584960 192628
rect 580901 192536 584960 192538
rect 580901 192480 580906 192536
rect 580962 192480 584960 192536
rect 580901 192478 584960 192480
rect 580901 192475 580967 192478
rect 583520 192388 584960 192478
rect 1301 192130 1367 192133
rect 1301 192128 3220 192130
rect 1301 192072 1306 192128
rect 1362 192072 3220 192128
rect 1301 192070 3220 192072
rect 1301 192067 1367 192070
rect -960 188866 480 188956
rect 1301 188866 1367 188869
rect -960 188864 1367 188866
rect -960 188808 1306 188864
rect 1362 188808 1367 188864
rect -960 188806 1367 188808
rect -960 188716 480 188806
rect 1301 188803 1367 188806
rect 580901 182474 580967 182477
rect 580766 182472 580967 182474
rect 580766 182416 580906 182472
rect 580962 182416 580967 182472
rect 580766 182414 580967 182416
rect 580766 182308 580826 182414
rect 580901 182411 580967 182414
rect 2773 179346 2839 179349
rect 2773 179344 3220 179346
rect 2773 179288 2778 179344
rect 2834 179288 3220 179344
rect 2773 179286 3220 179288
rect 2773 179283 2839 179286
rect 580901 179210 580967 179213
rect 583520 179210 584960 179300
rect 580901 179208 584960 179210
rect 580901 179152 580906 179208
rect 580962 179152 584960 179208
rect 580901 179150 584960 179152
rect 580901 179147 580967 179150
rect 583520 179060 584960 179150
rect -960 175946 480 176036
rect 2773 175946 2839 175949
rect -960 175944 2839 175946
rect -960 175888 2778 175944
rect 2834 175888 2839 175944
rect -960 175886 2839 175888
rect -960 175796 480 175886
rect 2773 175883 2839 175886
rect 580766 168602 580826 169116
rect 580901 168602 580967 168605
rect 580766 168600 580967 168602
rect 580766 168544 580906 168600
rect 580962 168544 580967 168600
rect 580766 168542 580967 168544
rect 580901 168539 580967 168542
rect 2773 166562 2839 166565
rect 2773 166560 3220 166562
rect 2773 166504 2778 166560
rect 2834 166504 3220 166560
rect 2773 166502 3220 166504
rect 2773 166499 2839 166502
rect 580901 165882 580967 165885
rect 583520 165882 584960 165972
rect 580901 165880 584960 165882
rect 580901 165824 580906 165880
rect 580962 165824 584960 165880
rect 580901 165822 584960 165824
rect 580901 165819 580967 165822
rect 583520 165732 584960 165822
rect -960 162890 480 162980
rect 2773 162890 2839 162893
rect -960 162888 2839 162890
rect -960 162832 2778 162888
rect 2834 162832 2839 162888
rect -960 162830 2839 162832
rect -960 162740 480 162830
rect 2773 162827 2839 162830
rect 580901 156362 580967 156365
rect 580766 156360 580967 156362
rect 580766 156304 580906 156360
rect 580962 156304 580967 156360
rect 580766 156302 580967 156304
rect 580766 156196 580826 156302
rect 580901 156299 580967 156302
rect 1301 153778 1367 153781
rect 1301 153776 3220 153778
rect 1301 153720 1306 153776
rect 1362 153720 3220 153776
rect 1301 153718 3220 153720
rect 1301 153715 1367 153718
rect 580901 152690 580967 152693
rect 583520 152690 584960 152780
rect 580901 152688 584960 152690
rect 580901 152632 580906 152688
rect 580962 152632 584960 152688
rect 580901 152630 584960 152632
rect 580901 152627 580967 152630
rect 583520 152540 584960 152630
rect -960 149834 480 149924
rect 1301 149834 1367 149837
rect -960 149832 1367 149834
rect -960 149776 1306 149832
rect 1362 149776 1367 149832
rect -960 149774 1367 149776
rect -960 149684 480 149774
rect 1301 149771 1367 149774
rect 580766 142626 580826 143004
rect 580901 142626 580967 142629
rect 580766 142624 580967 142626
rect 580766 142568 580906 142624
rect 580962 142568 580967 142624
rect 580766 142566 580967 142568
rect 580901 142563 580967 142566
rect 565 140994 631 140997
rect 565 140992 3220 140994
rect 565 140936 570 140992
rect 626 140936 3220 140992
rect 565 140934 3220 140936
rect 565 140931 631 140934
rect 580901 139362 580967 139365
rect 583520 139362 584960 139452
rect 580901 139360 584960 139362
rect 580901 139304 580906 139360
rect 580962 139304 584960 139360
rect 580901 139302 584960 139304
rect 580901 139299 580967 139302
rect 583520 139212 584960 139302
rect -960 136778 480 136868
rect 565 136778 631 136781
rect -960 136776 631 136778
rect -960 136720 570 136776
rect 626 136720 631 136776
rect -960 136718 631 136720
rect -960 136628 480 136718
rect 565 136715 631 136718
rect 580901 130250 580967 130253
rect 580766 130248 580967 130250
rect 580766 130192 580906 130248
rect 580962 130192 580967 130248
rect 580766 130190 580967 130192
rect 580766 130084 580826 130190
rect 580901 130187 580967 130190
rect 749 128210 815 128213
rect 749 128208 3220 128210
rect 749 128152 754 128208
rect 810 128152 3220 128208
rect 749 128150 3220 128152
rect 749 128147 815 128150
rect 580901 126034 580967 126037
rect 583520 126034 584960 126124
rect 580901 126032 584960 126034
rect 580901 125976 580906 126032
rect 580962 125976 584960 126032
rect 580901 125974 584960 125976
rect 580901 125971 580967 125974
rect 583520 125884 584960 125974
rect -960 123722 480 123812
rect 749 123722 815 123725
rect -960 123720 815 123722
rect -960 123664 754 123720
rect 810 123664 815 123720
rect -960 123662 815 123664
rect -960 123572 480 123662
rect 749 123659 815 123662
rect 579889 116378 579955 116381
rect 580030 116378 580090 116892
rect 579889 116376 580090 116378
rect 579889 116320 579894 116376
rect 579950 116320 580090 116376
rect 579889 116318 580090 116320
rect 579889 116315 579955 116318
rect 1301 115426 1367 115429
rect 1301 115424 3220 115426
rect 1301 115368 1306 115424
rect 1362 115368 3220 115424
rect 1301 115366 3220 115368
rect 1301 115363 1367 115366
rect 579889 112842 579955 112845
rect 583520 112842 584960 112932
rect 579889 112840 584960 112842
rect 579889 112784 579894 112840
rect 579950 112784 584960 112840
rect 579889 112782 584960 112784
rect 579889 112779 579955 112782
rect 583520 112692 584960 112782
rect -960 110666 480 110756
rect 1301 110666 1367 110669
rect -960 110664 1367 110666
rect -960 110608 1306 110664
rect 1362 110608 1367 110664
rect -960 110606 1367 110608
rect -960 110516 480 110606
rect 1301 110603 1367 110606
rect 580766 103594 580826 103836
rect 580901 103594 580967 103597
rect 580766 103592 580967 103594
rect 580766 103536 580906 103592
rect 580962 103536 580967 103592
rect 580766 103534 580967 103536
rect 580901 103531 580967 103534
rect 1577 102642 1643 102645
rect 1577 102640 3220 102642
rect 1577 102584 1582 102640
rect 1638 102584 3220 102640
rect 1577 102582 3220 102584
rect 1577 102579 1643 102582
rect 580901 99514 580967 99517
rect 583520 99514 584960 99604
rect 580901 99512 584960 99514
rect 580901 99456 580906 99512
rect 580962 99456 584960 99512
rect 580901 99454 584960 99456
rect 580901 99451 580967 99454
rect 583520 99364 584960 99454
rect -960 97610 480 97700
rect 1577 97610 1643 97613
rect -960 97608 1643 97610
rect -960 97552 1582 97608
rect 1638 97552 1643 97608
rect -960 97550 1643 97552
rect -960 97460 480 97550
rect 1577 97547 1643 97550
rect 580766 90266 580826 90780
rect 580901 90266 580967 90269
rect 580766 90264 580967 90266
rect 580766 90208 580906 90264
rect 580962 90208 580967 90264
rect 580766 90206 580967 90208
rect 580901 90203 580967 90206
rect 1577 89858 1643 89861
rect 1577 89856 3220 89858
rect 1577 89800 1582 89856
rect 1638 89800 3220 89856
rect 1577 89798 3220 89800
rect 1577 89795 1643 89798
rect 580901 86186 580967 86189
rect 583520 86186 584960 86276
rect 580901 86184 584960 86186
rect 580901 86128 580906 86184
rect 580962 86128 584960 86184
rect 580901 86126 584960 86128
rect 580901 86123 580967 86126
rect 583520 86036 584960 86126
rect -960 84690 480 84780
rect 1577 84690 1643 84693
rect -960 84688 1643 84690
rect -960 84632 1582 84688
rect 1638 84632 1643 84688
rect -960 84630 1643 84632
rect -960 84540 480 84630
rect 1577 84627 1643 84630
rect 579889 77346 579955 77349
rect 580030 77346 580090 77724
rect 579889 77344 580090 77346
rect 579889 77288 579894 77344
rect 579950 77288 580090 77344
rect 579889 77286 580090 77288
rect 579889 77283 579955 77286
rect 1577 77074 1643 77077
rect 1577 77072 3220 77074
rect 1577 77016 1582 77072
rect 1638 77016 3220 77072
rect 1577 77014 3220 77016
rect 1577 77011 1643 77014
rect 579889 72994 579955 72997
rect 583520 72994 584960 73084
rect 579889 72992 584960 72994
rect 579889 72936 579894 72992
rect 579950 72936 584960 72992
rect 579889 72934 584960 72936
rect 579889 72931 579955 72934
rect 583520 72844 584960 72934
rect -960 71634 480 71724
rect 1577 71634 1643 71637
rect -960 71632 1643 71634
rect -960 71576 1582 71632
rect 1638 71576 1643 71632
rect -960 71574 1643 71576
rect -960 71484 480 71574
rect 1577 71571 1643 71574
rect 1485 64290 1551 64293
rect 1485 64288 3220 64290
rect 1485 64232 1490 64288
rect 1546 64232 3220 64288
rect 1485 64230 3220 64232
rect 1485 64227 1551 64230
rect 580766 64154 580826 64668
rect 580901 64154 580967 64157
rect 580766 64152 580967 64154
rect 580766 64096 580906 64152
rect 580962 64096 580967 64152
rect 580766 64094 580967 64096
rect 580901 64091 580967 64094
rect 580901 59666 580967 59669
rect 583520 59666 584960 59756
rect 580901 59664 584960 59666
rect 580901 59608 580906 59664
rect 580962 59608 584960 59664
rect 580901 59606 584960 59608
rect 580901 59603 580967 59606
rect 583520 59516 584960 59606
rect -960 58578 480 58668
rect 1485 58578 1551 58581
rect -960 58576 1551 58578
rect -960 58520 1490 58576
rect 1546 58520 1551 58576
rect -960 58518 1551 58520
rect -960 58428 480 58518
rect 1485 58515 1551 58518
rect 2037 51506 2103 51509
rect 2037 51504 3220 51506
rect 2037 51448 2042 51504
rect 2098 51448 3220 51504
rect 2037 51446 3220 51448
rect 2037 51443 2103 51446
rect 580766 51098 580826 51612
rect 580901 51098 580967 51101
rect 580766 51096 580967 51098
rect 580766 51040 580906 51096
rect 580962 51040 580967 51096
rect 580766 51038 580967 51040
rect 580901 51035 580967 51038
rect 580901 46338 580967 46341
rect 583520 46338 584960 46428
rect 580901 46336 584960 46338
rect 580901 46280 580906 46336
rect 580962 46280 584960 46336
rect 580901 46278 584960 46280
rect 580901 46275 580967 46278
rect 583520 46188 584960 46278
rect -960 45522 480 45612
rect 2037 45522 2103 45525
rect -960 45520 2103 45522
rect -960 45464 2042 45520
rect 2098 45464 2103 45520
rect -960 45462 2103 45464
rect -960 45372 480 45462
rect 2037 45459 2103 45462
rect 2037 38722 2103 38725
rect 2037 38720 3220 38722
rect 2037 38664 2042 38720
rect 2098 38664 3220 38720
rect 2037 38662 3220 38664
rect 2037 38659 2103 38662
rect 580766 38042 580826 38556
rect 580901 38042 580967 38045
rect 580766 38040 580967 38042
rect 580766 37984 580906 38040
rect 580962 37984 580967 38040
rect 580766 37982 580967 37984
rect 580901 37979 580967 37982
rect 580901 33146 580967 33149
rect 583520 33146 584960 33236
rect 580901 33144 584960 33146
rect 580901 33088 580906 33144
rect 580962 33088 584960 33144
rect 580901 33086 584960 33088
rect 580901 33083 580967 33086
rect 583520 32996 584960 33086
rect -960 32466 480 32556
rect 2037 32466 2103 32469
rect -960 32464 2103 32466
rect -960 32408 2042 32464
rect 2098 32408 2103 32464
rect -960 32406 2103 32408
rect -960 32316 480 32406
rect 2037 32403 2103 32406
rect 1485 25938 1551 25941
rect 1485 25936 3220 25938
rect 1485 25880 1490 25936
rect 1546 25880 3220 25936
rect 1485 25878 3220 25880
rect 1485 25875 1551 25878
rect 580766 24986 580826 25500
rect 580901 24986 580967 24989
rect 580766 24984 580967 24986
rect 580766 24928 580906 24984
rect 580962 24928 580967 24984
rect 580766 24926 580967 24928
rect 580901 24923 580967 24926
rect 580901 19818 580967 19821
rect 583520 19818 584960 19908
rect 580901 19816 584960 19818
rect 580901 19760 580906 19816
rect 580962 19760 584960 19816
rect 580901 19758 584960 19760
rect 580901 19755 580967 19758
rect 583520 19668 584960 19758
rect -960 19410 480 19500
rect 1485 19410 1551 19413
rect -960 19408 1551 19410
rect -960 19352 1490 19408
rect 1546 19352 1551 19408
rect -960 19350 1551 19352
rect -960 19260 480 19350
rect 1485 19347 1551 19350
rect 2037 13154 2103 13157
rect 2037 13152 3220 13154
rect 2037 13096 2042 13152
rect 2098 13096 3220 13152
rect 2037 13094 3220 13096
rect 2037 13091 2103 13094
rect 579889 12746 579955 12749
rect 579889 12744 580090 12746
rect 579889 12688 579894 12744
rect 579950 12688 580090 12744
rect 579889 12686 580090 12688
rect 579889 12683 579955 12686
rect 580030 12580 580090 12686
rect 579889 6626 579955 6629
rect 583520 6626 584960 6716
rect 579889 6624 584960 6626
rect -960 6490 480 6580
rect 579889 6568 579894 6624
rect 579950 6568 584960 6624
rect 579889 6566 584960 6568
rect 579889 6563 579955 6566
rect 2037 6490 2103 6493
rect -960 6488 2103 6490
rect -960 6432 2042 6488
rect 2098 6432 2103 6488
rect 583520 6476 584960 6566
rect -960 6430 2103 6432
rect -960 6340 480 6430
rect 2037 6427 2103 6430
rect 70209 3906 70275 3909
rect 73613 3906 73679 3909
rect 70209 3904 73679 3906
rect 70209 3848 70214 3904
rect 70270 3848 73618 3904
rect 73674 3848 73679 3904
rect 70209 3846 73679 3848
rect 70209 3843 70275 3846
rect 73613 3843 73679 3846
rect 28901 642 28967 645
rect 46289 642 46355 645
rect 28901 640 46355 642
rect 28901 584 28906 640
rect 28962 584 46294 640
rect 46350 584 46355 640
rect 28901 582 46355 584
rect 28901 579 28967 582
rect 46289 579 46355 582
rect 12157 506 12223 509
rect 30833 506 30899 509
rect 12157 504 30899 506
rect 12157 448 12162 504
rect 12218 448 30838 504
rect 30894 448 30899 504
rect 12157 446 30899 448
rect 12157 443 12223 446
rect 30833 443 30899 446
rect 5441 370 5507 373
rect 23933 370 23999 373
rect 5441 368 23999 370
rect 5441 312 5446 368
rect 5502 312 23938 368
rect 23994 312 23999 368
rect 5441 310 23999 312
rect 5441 307 5507 310
rect 23933 307 23999 310
rect 25681 370 25747 373
rect 42701 370 42767 373
rect 25681 368 42767 370
rect 25681 312 25686 368
rect 25742 312 42706 368
rect 42762 312 42767 368
rect 25681 310 42767 312
rect 25681 307 25747 310
rect 42701 307 42767 310
rect 13721 234 13787 237
rect 31937 234 32003 237
rect 13721 232 32003 234
rect 13721 176 13726 232
rect 13782 176 31942 232
rect 31998 176 32003 232
rect 13721 174 32003 176
rect 13721 171 13787 174
rect 31937 171 32003 174
rect 36997 234 37063 237
rect 54017 234 54083 237
rect 36997 232 54083 234
rect 36997 176 37002 232
rect 37058 176 54022 232
rect 54078 176 54083 232
rect 36997 174 54083 176
rect 36997 171 37063 174
rect 54017 171 54083 174
rect 6269 98 6335 101
rect 25037 98 25103 101
rect 6269 96 25103 98
rect 6269 40 6274 96
rect 6330 40 25042 96
rect 25098 40 25103 96
rect 6269 38 25103 40
rect 6269 35 6335 38
rect 25037 35 25103 38
rect 46841 98 46907 101
rect 62849 98 62915 101
rect 46841 96 62915 98
rect 46841 40 46846 96
rect 46902 40 62854 96
rect 62910 40 62915 96
rect 46841 38 62915 40
rect 46841 35 46907 38
rect 62849 35 62915 38
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 -7066 -8106 711002
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 -6106 -7146 710042
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 -5146 -6186 709082
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 -4186 -5226 708122
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 -3226 -4266 707162
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 -2266 -3306 706202
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 700954 -2346 705242
rect 582294 705798 582914 711590
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 582294 705562 582326 705798
rect 582562 705562 582646 705798
rect 582882 705562 582914 705798
rect 582294 705478 582914 705562
rect 582294 705242 582326 705478
rect 582562 705242 582646 705478
rect 582882 705242 582914 705478
rect -2966 700718 -2934 700954
rect -2698 700718 -2614 700954
rect -2378 700718 -2346 700954
rect -2966 700634 -2346 700718
rect -2966 700398 -2934 700634
rect -2698 700398 -2614 700634
rect -2378 700398 -2346 700634
rect -2966 664954 -2346 700398
rect -2966 664718 -2934 664954
rect -2698 664718 -2614 664954
rect -2378 664718 -2346 664954
rect -2966 664634 -2346 664718
rect -2966 664398 -2934 664634
rect -2698 664398 -2614 664634
rect -2378 664398 -2346 664634
rect -2966 628954 -2346 664398
rect -2966 628718 -2934 628954
rect -2698 628718 -2614 628954
rect -2378 628718 -2346 628954
rect -2966 628634 -2346 628718
rect -2966 628398 -2934 628634
rect -2698 628398 -2614 628634
rect -2378 628398 -2346 628634
rect -2966 592954 -2346 628398
rect -2966 592718 -2934 592954
rect -2698 592718 -2614 592954
rect -2378 592718 -2346 592954
rect -2966 592634 -2346 592718
rect -2966 592398 -2934 592634
rect -2698 592398 -2614 592634
rect -2378 592398 -2346 592634
rect -2966 556954 -2346 592398
rect -2966 556718 -2934 556954
rect -2698 556718 -2614 556954
rect -2378 556718 -2346 556954
rect -2966 556634 -2346 556718
rect -2966 556398 -2934 556634
rect -2698 556398 -2614 556634
rect -2378 556398 -2346 556634
rect -2966 520954 -2346 556398
rect -2966 520718 -2934 520954
rect -2698 520718 -2614 520954
rect -2378 520718 -2346 520954
rect -2966 520634 -2346 520718
rect -2966 520398 -2934 520634
rect -2698 520398 -2614 520634
rect -2378 520398 -2346 520634
rect -2966 484954 -2346 520398
rect -2966 484718 -2934 484954
rect -2698 484718 -2614 484954
rect -2378 484718 -2346 484954
rect -2966 484634 -2346 484718
rect -2966 484398 -2934 484634
rect -2698 484398 -2614 484634
rect -2378 484398 -2346 484634
rect -2966 448954 -2346 484398
rect -2966 448718 -2934 448954
rect -2698 448718 -2614 448954
rect -2378 448718 -2346 448954
rect -2966 448634 -2346 448718
rect -2966 448398 -2934 448634
rect -2698 448398 -2614 448634
rect -2378 448398 -2346 448634
rect -2966 412954 -2346 448398
rect -2966 412718 -2934 412954
rect -2698 412718 -2614 412954
rect -2378 412718 -2346 412954
rect -2966 412634 -2346 412718
rect -2966 412398 -2934 412634
rect -2698 412398 -2614 412634
rect -2378 412398 -2346 412634
rect -2966 376954 -2346 412398
rect -2966 376718 -2934 376954
rect -2698 376718 -2614 376954
rect -2378 376718 -2346 376954
rect -2966 376634 -2346 376718
rect -2966 376398 -2934 376634
rect -2698 376398 -2614 376634
rect -2378 376398 -2346 376634
rect -2966 340954 -2346 376398
rect -2966 340718 -2934 340954
rect -2698 340718 -2614 340954
rect -2378 340718 -2346 340954
rect -2966 340634 -2346 340718
rect -2966 340398 -2934 340634
rect -2698 340398 -2614 340634
rect -2378 340398 -2346 340634
rect -2966 304954 -2346 340398
rect -2966 304718 -2934 304954
rect -2698 304718 -2614 304954
rect -2378 304718 -2346 304954
rect -2966 304634 -2346 304718
rect -2966 304398 -2934 304634
rect -2698 304398 -2614 304634
rect -2378 304398 -2346 304634
rect -2966 268954 -2346 304398
rect -2966 268718 -2934 268954
rect -2698 268718 -2614 268954
rect -2378 268718 -2346 268954
rect -2966 268634 -2346 268718
rect -2966 268398 -2934 268634
rect -2698 268398 -2614 268634
rect -2378 268398 -2346 268634
rect -2966 232954 -2346 268398
rect -2966 232718 -2934 232954
rect -2698 232718 -2614 232954
rect -2378 232718 -2346 232954
rect -2966 232634 -2346 232718
rect -2966 232398 -2934 232634
rect -2698 232398 -2614 232634
rect -2378 232398 -2346 232634
rect -2966 196954 -2346 232398
rect -2966 196718 -2934 196954
rect -2698 196718 -2614 196954
rect -2378 196718 -2346 196954
rect -2966 196634 -2346 196718
rect -2966 196398 -2934 196634
rect -2698 196398 -2614 196634
rect -2378 196398 -2346 196634
rect -2966 160954 -2346 196398
rect -2966 160718 -2934 160954
rect -2698 160718 -2614 160954
rect -2378 160718 -2346 160954
rect -2966 160634 -2346 160718
rect -2966 160398 -2934 160634
rect -2698 160398 -2614 160634
rect -2378 160398 -2346 160634
rect -2966 124954 -2346 160398
rect -2966 124718 -2934 124954
rect -2698 124718 -2614 124954
rect -2378 124718 -2346 124954
rect -2966 124634 -2346 124718
rect -2966 124398 -2934 124634
rect -2698 124398 -2614 124634
rect -2378 124398 -2346 124634
rect -2966 88954 -2346 124398
rect -2966 88718 -2934 88954
rect -2698 88718 -2614 88954
rect -2378 88718 -2346 88954
rect -2966 88634 -2346 88718
rect -2966 88398 -2934 88634
rect -2698 88398 -2614 88634
rect -2378 88398 -2346 88634
rect -2966 52954 -2346 88398
rect -2966 52718 -2934 52954
rect -2698 52718 -2614 52954
rect -2378 52718 -2346 52954
rect -2966 52634 -2346 52718
rect -2966 52398 -2934 52634
rect -2698 52398 -2614 52634
rect -2378 52398 -2346 52634
rect -2966 16954 -2346 52398
rect -2966 16718 -2934 16954
rect -2698 16718 -2614 16954
rect -2378 16718 -2346 16954
rect -2966 16634 -2346 16718
rect -2966 16398 -2934 16634
rect -2698 16398 -2614 16634
rect -2378 16398 -2346 16634
rect -2966 -1306 -2346 16398
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 696454 -1386 704282
rect 582294 700954 582914 705242
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 582294 700718 582326 700954
rect 582562 700718 582646 700954
rect 582882 700718 582914 700954
rect 582294 700634 582914 700718
rect 582294 700398 582326 700634
rect 582562 700398 582646 700634
rect 582882 700398 582914 700634
rect -2006 696218 -1974 696454
rect -1738 696218 -1654 696454
rect -1418 696218 -1386 696454
rect -2006 696134 -1386 696218
rect -2006 695898 -1974 696134
rect -1738 695898 -1654 696134
rect -1418 695898 -1386 696134
rect 5794 696218 5826 696454
rect 6062 696218 6146 696454
rect 6382 696218 6414 696454
rect 5794 696134 6414 696218
rect 5794 695898 5826 696134
rect 6062 695898 6146 696134
rect 6382 695898 6414 696134
rect 41794 696218 41826 696454
rect 42062 696218 42146 696454
rect 42382 696218 42414 696454
rect 41794 696134 42414 696218
rect 41794 695898 41826 696134
rect 42062 695898 42146 696134
rect 42382 695898 42414 696134
rect 77794 696218 77826 696454
rect 78062 696218 78146 696454
rect 78382 696218 78414 696454
rect 77794 696134 78414 696218
rect 77794 695898 77826 696134
rect 78062 695898 78146 696134
rect 78382 695898 78414 696134
rect 113794 696218 113826 696454
rect 114062 696218 114146 696454
rect 114382 696218 114414 696454
rect 113794 696134 114414 696218
rect 113794 695898 113826 696134
rect 114062 695898 114146 696134
rect 114382 695898 114414 696134
rect 149794 696218 149826 696454
rect 150062 696218 150146 696454
rect 150382 696218 150414 696454
rect 149794 696134 150414 696218
rect 149794 695898 149826 696134
rect 150062 695898 150146 696134
rect 150382 695898 150414 696134
rect 185794 696218 185826 696454
rect 186062 696218 186146 696454
rect 186382 696218 186414 696454
rect 185794 696134 186414 696218
rect 185794 695898 185826 696134
rect 186062 695898 186146 696134
rect 186382 695898 186414 696134
rect 221794 696218 221826 696454
rect 222062 696218 222146 696454
rect 222382 696218 222414 696454
rect 221794 696134 222414 696218
rect 221794 695898 221826 696134
rect 222062 695898 222146 696134
rect 222382 695898 222414 696134
rect 257794 696218 257826 696454
rect 258062 696218 258146 696454
rect 258382 696218 258414 696454
rect 257794 696134 258414 696218
rect 257794 695898 257826 696134
rect 258062 695898 258146 696134
rect 258382 695898 258414 696134
rect 293794 696218 293826 696454
rect 294062 696218 294146 696454
rect 294382 696218 294414 696454
rect 293794 696134 294414 696218
rect 293794 695898 293826 696134
rect 294062 695898 294146 696134
rect 294382 695898 294414 696134
rect 329794 696218 329826 696454
rect 330062 696218 330146 696454
rect 330382 696218 330414 696454
rect 329794 696134 330414 696218
rect 329794 695898 329826 696134
rect 330062 695898 330146 696134
rect 330382 695898 330414 696134
rect 365794 696218 365826 696454
rect 366062 696218 366146 696454
rect 366382 696218 366414 696454
rect 365794 696134 366414 696218
rect 365794 695898 365826 696134
rect 366062 695898 366146 696134
rect 366382 695898 366414 696134
rect 401794 696218 401826 696454
rect 402062 696218 402146 696454
rect 402382 696218 402414 696454
rect 401794 696134 402414 696218
rect 401794 695898 401826 696134
rect 402062 695898 402146 696134
rect 402382 695898 402414 696134
rect 437794 696218 437826 696454
rect 438062 696218 438146 696454
rect 438382 696218 438414 696454
rect 437794 696134 438414 696218
rect 437794 695898 437826 696134
rect 438062 695898 438146 696134
rect 438382 695898 438414 696134
rect 473794 696218 473826 696454
rect 474062 696218 474146 696454
rect 474382 696218 474414 696454
rect 473794 696134 474414 696218
rect 473794 695898 473826 696134
rect 474062 695898 474146 696134
rect 474382 695898 474414 696134
rect 509794 696218 509826 696454
rect 510062 696218 510146 696454
rect 510382 696218 510414 696454
rect 509794 696134 510414 696218
rect 509794 695898 509826 696134
rect 510062 695898 510146 696134
rect 510382 695898 510414 696134
rect 545794 696218 545826 696454
rect 546062 696218 546146 696454
rect 546382 696218 546414 696454
rect 545794 696134 546414 696218
rect 545794 695898 545826 696134
rect 546062 695898 546146 696134
rect 546382 695898 546414 696134
rect -2006 660454 -1386 695898
rect 582294 664954 582914 700398
rect 13166 664718 13198 664954
rect 13434 664718 13518 664954
rect 13754 664718 13786 664954
rect 13166 664634 13786 664718
rect 13166 664398 13198 664634
rect 13434 664398 13518 664634
rect 13754 664398 13786 664634
rect 167794 664718 167826 664954
rect 168062 664718 168146 664954
rect 168382 664718 168414 664954
rect 167794 664634 168414 664718
rect 167794 664398 167826 664634
rect 168062 664398 168146 664634
rect 168382 664398 168414 664634
rect 291558 664718 291590 664954
rect 291826 664718 291910 664954
rect 292146 664718 292178 664954
rect 291558 664634 292178 664718
rect 291558 664398 291590 664634
rect 291826 664398 291910 664634
rect 292146 664398 292178 664634
rect 419794 664718 419826 664954
rect 420062 664718 420146 664954
rect 420382 664718 420414 664954
rect 419794 664634 420414 664718
rect 419794 664398 419826 664634
rect 420062 664398 420146 664634
rect 420382 664398 420414 664634
rect 563794 664718 563826 664954
rect 564062 664718 564146 664954
rect 564382 664718 564414 664954
rect 563794 664634 564414 664718
rect 563794 664398 563826 664634
rect 564062 664398 564146 664634
rect 564382 664398 564414 664634
rect 582294 664718 582326 664954
rect 582562 664718 582646 664954
rect 582882 664718 582914 664954
rect 582294 664634 582914 664718
rect 582294 664398 582326 664634
rect 582562 664398 582646 664634
rect 582882 664398 582914 664634
rect -2006 660218 -1974 660454
rect -1738 660218 -1654 660454
rect -1418 660218 -1386 660454
rect -2006 660134 -1386 660218
rect -2006 659898 -1974 660134
rect -1738 659898 -1654 660134
rect -1418 659898 -1386 660134
rect 5794 660218 5826 660454
rect 6062 660218 6146 660454
rect 6382 660218 6414 660454
rect 5794 660134 6414 660218
rect 5794 659898 5826 660134
rect 6062 659898 6146 660134
rect 6382 659898 6414 660134
rect 173062 660218 173094 660454
rect 173330 660218 173414 660454
rect 173650 660218 173682 660454
rect 173062 660134 173682 660218
rect 173062 659898 173094 660134
rect 173330 659898 173414 660134
rect 173650 659898 173682 660134
rect 293794 660218 293826 660454
rect 294062 660218 294146 660454
rect 294382 660218 294414 660454
rect 293794 660134 294414 660218
rect 293794 659898 293826 660134
rect 294062 659898 294146 660134
rect 294382 659898 294414 660134
rect 401794 660218 401826 660454
rect 402062 660218 402146 660454
rect 402382 660218 402414 660454
rect 401794 660134 402414 660218
rect 401794 659898 401826 660134
rect 402062 659898 402146 660134
rect 402382 659898 402414 660134
rect 570318 660218 570350 660454
rect 570586 660218 570670 660454
rect 570906 660218 570938 660454
rect 570318 660134 570938 660218
rect 570318 659898 570350 660134
rect 570586 659898 570670 660134
rect 570906 659898 570938 660134
rect -2006 624454 -1386 659898
rect 582294 628954 582914 664398
rect 13166 628718 13198 628954
rect 13434 628718 13518 628954
rect 13754 628718 13786 628954
rect 13166 628634 13786 628718
rect 13166 628398 13198 628634
rect 13434 628398 13518 628634
rect 13754 628398 13786 628634
rect 167794 628718 167826 628954
rect 168062 628718 168146 628954
rect 168382 628718 168414 628954
rect 167794 628634 168414 628718
rect 167794 628398 167826 628634
rect 168062 628398 168146 628634
rect 168382 628398 168414 628634
rect 291558 628718 291590 628954
rect 291826 628718 291910 628954
rect 292146 628718 292178 628954
rect 291558 628634 292178 628718
rect 291558 628398 291590 628634
rect 291826 628398 291910 628634
rect 292146 628398 292178 628634
rect 419794 628718 419826 628954
rect 420062 628718 420146 628954
rect 420382 628718 420414 628954
rect 419794 628634 420414 628718
rect 419794 628398 419826 628634
rect 420062 628398 420146 628634
rect 420382 628398 420414 628634
rect 563794 628718 563826 628954
rect 564062 628718 564146 628954
rect 564382 628718 564414 628954
rect 563794 628634 564414 628718
rect 563794 628398 563826 628634
rect 564062 628398 564146 628634
rect 564382 628398 564414 628634
rect 582294 628718 582326 628954
rect 582562 628718 582646 628954
rect 582882 628718 582914 628954
rect 582294 628634 582914 628718
rect 582294 628398 582326 628634
rect 582562 628398 582646 628634
rect 582882 628398 582914 628634
rect -2006 624218 -1974 624454
rect -1738 624218 -1654 624454
rect -1418 624218 -1386 624454
rect -2006 624134 -1386 624218
rect -2006 623898 -1974 624134
rect -1738 623898 -1654 624134
rect -1418 623898 -1386 624134
rect 5794 624218 5826 624454
rect 6062 624218 6146 624454
rect 6382 624218 6414 624454
rect 5794 624134 6414 624218
rect 5794 623898 5826 624134
rect 6062 623898 6146 624134
rect 6382 623898 6414 624134
rect 173062 624218 173094 624454
rect 173330 624218 173414 624454
rect 173650 624218 173682 624454
rect 173062 624134 173682 624218
rect 173062 623898 173094 624134
rect 173330 623898 173414 624134
rect 173650 623898 173682 624134
rect 293794 624218 293826 624454
rect 294062 624218 294146 624454
rect 294382 624218 294414 624454
rect 293794 624134 294414 624218
rect 293794 623898 293826 624134
rect 294062 623898 294146 624134
rect 294382 623898 294414 624134
rect 401794 624218 401826 624454
rect 402062 624218 402146 624454
rect 402382 624218 402414 624454
rect 401794 624134 402414 624218
rect 401794 623898 401826 624134
rect 402062 623898 402146 624134
rect 402382 623898 402414 624134
rect 570318 624218 570350 624454
rect 570586 624218 570670 624454
rect 570906 624218 570938 624454
rect 570318 624134 570938 624218
rect 570318 623898 570350 624134
rect 570586 623898 570670 624134
rect 570906 623898 570938 624134
rect -2006 588454 -1386 623898
rect 582294 592954 582914 628398
rect 23794 592718 23826 592954
rect 24062 592718 24146 592954
rect 24382 592718 24414 592954
rect 23794 592634 24414 592718
rect 23794 592398 23826 592634
rect 24062 592398 24146 592634
rect 24382 592398 24414 592634
rect 59794 592718 59826 592954
rect 60062 592718 60146 592954
rect 60382 592718 60414 592954
rect 59794 592634 60414 592718
rect 59794 592398 59826 592634
rect 60062 592398 60146 592634
rect 60382 592398 60414 592634
rect 95794 592718 95826 592954
rect 96062 592718 96146 592954
rect 96382 592718 96414 592954
rect 95794 592634 96414 592718
rect 95794 592398 95826 592634
rect 96062 592398 96146 592634
rect 96382 592398 96414 592634
rect 131794 592718 131826 592954
rect 132062 592718 132146 592954
rect 132382 592718 132414 592954
rect 131794 592634 132414 592718
rect 131794 592398 131826 592634
rect 132062 592398 132146 592634
rect 132382 592398 132414 592634
rect 167794 592718 167826 592954
rect 168062 592718 168146 592954
rect 168382 592718 168414 592954
rect 167794 592634 168414 592718
rect 167794 592398 167826 592634
rect 168062 592398 168146 592634
rect 168382 592398 168414 592634
rect 291558 592718 291590 592954
rect 291826 592718 291910 592954
rect 292146 592718 292178 592954
rect 291558 592634 292178 592718
rect 291558 592398 291590 592634
rect 291826 592398 291910 592634
rect 292146 592398 292178 592634
rect 419794 592718 419826 592954
rect 420062 592718 420146 592954
rect 420382 592718 420414 592954
rect 419794 592634 420414 592718
rect 419794 592398 419826 592634
rect 420062 592398 420146 592634
rect 420382 592398 420414 592634
rect 455794 592718 455826 592954
rect 456062 592718 456146 592954
rect 456382 592718 456414 592954
rect 455794 592634 456414 592718
rect 455794 592398 455826 592634
rect 456062 592398 456146 592634
rect 456382 592398 456414 592634
rect 491794 592718 491826 592954
rect 492062 592718 492146 592954
rect 492382 592718 492414 592954
rect 491794 592634 492414 592718
rect 491794 592398 491826 592634
rect 492062 592398 492146 592634
rect 492382 592398 492414 592634
rect 527794 592718 527826 592954
rect 528062 592718 528146 592954
rect 528382 592718 528414 592954
rect 527794 592634 528414 592718
rect 527794 592398 527826 592634
rect 528062 592398 528146 592634
rect 528382 592398 528414 592634
rect 563794 592718 563826 592954
rect 564062 592718 564146 592954
rect 564382 592718 564414 592954
rect 563794 592634 564414 592718
rect 563794 592398 563826 592634
rect 564062 592398 564146 592634
rect 564382 592398 564414 592634
rect 582294 592718 582326 592954
rect 582562 592718 582646 592954
rect 582882 592718 582914 592954
rect 582294 592634 582914 592718
rect 582294 592398 582326 592634
rect 582562 592398 582646 592634
rect 582882 592398 582914 592634
rect -2006 588218 -1974 588454
rect -1738 588218 -1654 588454
rect -1418 588218 -1386 588454
rect -2006 588134 -1386 588218
rect -2006 587898 -1974 588134
rect -1738 587898 -1654 588134
rect -1418 587898 -1386 588134
rect 5794 588218 5826 588454
rect 6062 588218 6146 588454
rect 6382 588218 6414 588454
rect 5794 588134 6414 588218
rect 5794 587898 5826 588134
rect 6062 587898 6146 588134
rect 6382 587898 6414 588134
rect 41794 588218 41826 588454
rect 42062 588218 42146 588454
rect 42382 588218 42414 588454
rect 41794 588134 42414 588218
rect 41794 587898 41826 588134
rect 42062 587898 42146 588134
rect 42382 587898 42414 588134
rect 77794 588218 77826 588454
rect 78062 588218 78146 588454
rect 78382 588218 78414 588454
rect 77794 588134 78414 588218
rect 77794 587898 77826 588134
rect 78062 587898 78146 588134
rect 78382 587898 78414 588134
rect 113794 588218 113826 588454
rect 114062 588218 114146 588454
rect 114382 588218 114414 588454
rect 113794 588134 114414 588218
rect 113794 587898 113826 588134
rect 114062 587898 114146 588134
rect 114382 587898 114414 588134
rect 149794 588218 149826 588454
rect 150062 588218 150146 588454
rect 150382 588218 150414 588454
rect 149794 588134 150414 588218
rect 149794 587898 149826 588134
rect 150062 587898 150146 588134
rect 150382 587898 150414 588134
rect 185794 588218 185826 588454
rect 186062 588218 186146 588454
rect 186382 588218 186414 588454
rect 185794 588134 186414 588218
rect 185794 587898 185826 588134
rect 186062 587898 186146 588134
rect 186382 587898 186414 588134
rect 221794 588218 221826 588454
rect 222062 588218 222146 588454
rect 222382 588218 222414 588454
rect 221794 588134 222414 588218
rect 221794 587898 221826 588134
rect 222062 587898 222146 588134
rect 222382 587898 222414 588134
rect 257794 588218 257826 588454
rect 258062 588218 258146 588454
rect 258382 588218 258414 588454
rect 257794 588134 258414 588218
rect 257794 587898 257826 588134
rect 258062 587898 258146 588134
rect 258382 587898 258414 588134
rect 293794 588218 293826 588454
rect 294062 588218 294146 588454
rect 294382 588218 294414 588454
rect 293794 588134 294414 588218
rect 293794 587898 293826 588134
rect 294062 587898 294146 588134
rect 294382 587898 294414 588134
rect 329794 588218 329826 588454
rect 330062 588218 330146 588454
rect 330382 588218 330414 588454
rect 329794 588134 330414 588218
rect 329794 587898 329826 588134
rect 330062 587898 330146 588134
rect 330382 587898 330414 588134
rect 365794 588218 365826 588454
rect 366062 588218 366146 588454
rect 366382 588218 366414 588454
rect 365794 588134 366414 588218
rect 365794 587898 365826 588134
rect 366062 587898 366146 588134
rect 366382 587898 366414 588134
rect 401794 588218 401826 588454
rect 402062 588218 402146 588454
rect 402382 588218 402414 588454
rect 401794 588134 402414 588218
rect 401794 587898 401826 588134
rect 402062 587898 402146 588134
rect 402382 587898 402414 588134
rect 437794 588218 437826 588454
rect 438062 588218 438146 588454
rect 438382 588218 438414 588454
rect 437794 588134 438414 588218
rect 437794 587898 437826 588134
rect 438062 587898 438146 588134
rect 438382 587898 438414 588134
rect 473794 588218 473826 588454
rect 474062 588218 474146 588454
rect 474382 588218 474414 588454
rect 473794 588134 474414 588218
rect 473794 587898 473826 588134
rect 474062 587898 474146 588134
rect 474382 587898 474414 588134
rect 509794 588218 509826 588454
rect 510062 588218 510146 588454
rect 510382 588218 510414 588454
rect 509794 588134 510414 588218
rect 509794 587898 509826 588134
rect 510062 587898 510146 588134
rect 510382 587898 510414 588134
rect 545794 588218 545826 588454
rect 546062 588218 546146 588454
rect 546382 588218 546414 588454
rect 545794 588134 546414 588218
rect 545794 587898 545826 588134
rect 546062 587898 546146 588134
rect 546382 587898 546414 588134
rect -2006 552454 -1386 587898
rect 582294 556954 582914 592398
rect 13166 556718 13198 556954
rect 13434 556718 13518 556954
rect 13754 556718 13786 556954
rect 13166 556634 13786 556718
rect 13166 556398 13198 556634
rect 13434 556398 13518 556634
rect 13754 556398 13786 556634
rect 167794 556718 167826 556954
rect 168062 556718 168146 556954
rect 168382 556718 168414 556954
rect 167794 556634 168414 556718
rect 167794 556398 167826 556634
rect 168062 556398 168146 556634
rect 168382 556398 168414 556634
rect 203794 556718 203826 556954
rect 204062 556718 204146 556954
rect 204382 556718 204414 556954
rect 203794 556634 204414 556718
rect 203794 556398 203826 556634
rect 204062 556398 204146 556634
rect 204382 556398 204414 556634
rect 239794 556718 239826 556954
rect 240062 556718 240146 556954
rect 240382 556718 240414 556954
rect 239794 556634 240414 556718
rect 239794 556398 239826 556634
rect 240062 556398 240146 556634
rect 240382 556398 240414 556634
rect 275794 556718 275826 556954
rect 276062 556718 276146 556954
rect 276382 556718 276414 556954
rect 275794 556634 276414 556718
rect 275794 556398 275826 556634
rect 276062 556398 276146 556634
rect 276382 556398 276414 556634
rect 311794 556718 311826 556954
rect 312062 556718 312146 556954
rect 312382 556718 312414 556954
rect 311794 556634 312414 556718
rect 311794 556398 311826 556634
rect 312062 556398 312146 556634
rect 312382 556398 312414 556634
rect 347794 556718 347826 556954
rect 348062 556718 348146 556954
rect 348382 556718 348414 556954
rect 347794 556634 348414 556718
rect 347794 556398 347826 556634
rect 348062 556398 348146 556634
rect 348382 556398 348414 556634
rect 383794 556718 383826 556954
rect 384062 556718 384146 556954
rect 384382 556718 384414 556954
rect 383794 556634 384414 556718
rect 383794 556398 383826 556634
rect 384062 556398 384146 556634
rect 384382 556398 384414 556634
rect 419794 556718 419826 556954
rect 420062 556718 420146 556954
rect 420382 556718 420414 556954
rect 419794 556634 420414 556718
rect 419794 556398 419826 556634
rect 420062 556398 420146 556634
rect 420382 556398 420414 556634
rect 563794 556718 563826 556954
rect 564062 556718 564146 556954
rect 564382 556718 564414 556954
rect 563794 556634 564414 556718
rect 563794 556398 563826 556634
rect 564062 556398 564146 556634
rect 564382 556398 564414 556634
rect 582294 556718 582326 556954
rect 582562 556718 582646 556954
rect 582882 556718 582914 556954
rect 582294 556634 582914 556718
rect 582294 556398 582326 556634
rect 582562 556398 582646 556634
rect 582882 556398 582914 556634
rect -2006 552218 -1974 552454
rect -1738 552218 -1654 552454
rect -1418 552218 -1386 552454
rect -2006 552134 -1386 552218
rect -2006 551898 -1974 552134
rect -1738 551898 -1654 552134
rect -1418 551898 -1386 552134
rect 5794 552218 5826 552454
rect 6062 552218 6146 552454
rect 6382 552218 6414 552454
rect 5794 552134 6414 552218
rect 5794 551898 5826 552134
rect 6062 551898 6146 552134
rect 6382 551898 6414 552134
rect 185794 552218 185826 552454
rect 186062 552218 186146 552454
rect 186382 552218 186414 552454
rect 185794 552134 186414 552218
rect 185794 551898 185826 552134
rect 186062 551898 186146 552134
rect 186382 551898 186414 552134
rect 221794 552218 221826 552454
rect 222062 552218 222146 552454
rect 222382 552218 222414 552454
rect 221794 552134 222414 552218
rect 221794 551898 221826 552134
rect 222062 551898 222146 552134
rect 222382 551898 222414 552134
rect 257794 552218 257826 552454
rect 258062 552218 258146 552454
rect 258382 552218 258414 552454
rect 257794 552134 258414 552218
rect 257794 551898 257826 552134
rect 258062 551898 258146 552134
rect 258382 551898 258414 552134
rect 293794 552218 293826 552454
rect 294062 552218 294146 552454
rect 294382 552218 294414 552454
rect 293794 552134 294414 552218
rect 293794 551898 293826 552134
rect 294062 551898 294146 552134
rect 294382 551898 294414 552134
rect 329794 552218 329826 552454
rect 330062 552218 330146 552454
rect 330382 552218 330414 552454
rect 329794 552134 330414 552218
rect 329794 551898 329826 552134
rect 330062 551898 330146 552134
rect 330382 551898 330414 552134
rect 365794 552218 365826 552454
rect 366062 552218 366146 552454
rect 366382 552218 366414 552454
rect 365794 552134 366414 552218
rect 365794 551898 365826 552134
rect 366062 551898 366146 552134
rect 366382 551898 366414 552134
rect 401794 552218 401826 552454
rect 402062 552218 402146 552454
rect 402382 552218 402414 552454
rect 401794 552134 402414 552218
rect 401794 551898 401826 552134
rect 402062 551898 402146 552134
rect 402382 551898 402414 552134
rect 570318 552218 570350 552454
rect 570586 552218 570670 552454
rect 570906 552218 570938 552454
rect 570318 552134 570938 552218
rect 570318 551898 570350 552134
rect 570586 551898 570670 552134
rect 570906 551898 570938 552134
rect -2006 516454 -1386 551898
rect 582294 520954 582914 556398
rect 13166 520718 13198 520954
rect 13434 520718 13518 520954
rect 13754 520718 13786 520954
rect 13166 520634 13786 520718
rect 13166 520398 13198 520634
rect 13434 520398 13518 520634
rect 13754 520398 13786 520634
rect 167794 520718 167826 520954
rect 168062 520718 168146 520954
rect 168382 520718 168414 520954
rect 167794 520634 168414 520718
rect 167794 520398 167826 520634
rect 168062 520398 168146 520634
rect 168382 520398 168414 520634
rect 203794 520718 203826 520954
rect 204062 520718 204146 520954
rect 204382 520718 204414 520954
rect 203794 520634 204414 520718
rect 203794 520398 203826 520634
rect 204062 520398 204146 520634
rect 204382 520398 204414 520634
rect 239794 520718 239826 520954
rect 240062 520718 240146 520954
rect 240382 520718 240414 520954
rect 239794 520634 240414 520718
rect 239794 520398 239826 520634
rect 240062 520398 240146 520634
rect 240382 520398 240414 520634
rect 275794 520718 275826 520954
rect 276062 520718 276146 520954
rect 276382 520718 276414 520954
rect 275794 520634 276414 520718
rect 275794 520398 275826 520634
rect 276062 520398 276146 520634
rect 276382 520398 276414 520634
rect 311794 520718 311826 520954
rect 312062 520718 312146 520954
rect 312382 520718 312414 520954
rect 311794 520634 312414 520718
rect 311794 520398 311826 520634
rect 312062 520398 312146 520634
rect 312382 520398 312414 520634
rect 347794 520718 347826 520954
rect 348062 520718 348146 520954
rect 348382 520718 348414 520954
rect 347794 520634 348414 520718
rect 347794 520398 347826 520634
rect 348062 520398 348146 520634
rect 348382 520398 348414 520634
rect 383794 520718 383826 520954
rect 384062 520718 384146 520954
rect 384382 520718 384414 520954
rect 383794 520634 384414 520718
rect 383794 520398 383826 520634
rect 384062 520398 384146 520634
rect 384382 520398 384414 520634
rect 419794 520718 419826 520954
rect 420062 520718 420146 520954
rect 420382 520718 420414 520954
rect 419794 520634 420414 520718
rect 419794 520398 419826 520634
rect 420062 520398 420146 520634
rect 420382 520398 420414 520634
rect 563794 520718 563826 520954
rect 564062 520718 564146 520954
rect 564382 520718 564414 520954
rect 563794 520634 564414 520718
rect 563794 520398 563826 520634
rect 564062 520398 564146 520634
rect 564382 520398 564414 520634
rect 582294 520718 582326 520954
rect 582562 520718 582646 520954
rect 582882 520718 582914 520954
rect 582294 520634 582914 520718
rect 582294 520398 582326 520634
rect 582562 520398 582646 520634
rect 582882 520398 582914 520634
rect -2006 516218 -1974 516454
rect -1738 516218 -1654 516454
rect -1418 516218 -1386 516454
rect -2006 516134 -1386 516218
rect -2006 515898 -1974 516134
rect -1738 515898 -1654 516134
rect -1418 515898 -1386 516134
rect 5794 516218 5826 516454
rect 6062 516218 6146 516454
rect 6382 516218 6414 516454
rect 5794 516134 6414 516218
rect 5794 515898 5826 516134
rect 6062 515898 6146 516134
rect 6382 515898 6414 516134
rect 185794 516218 185826 516454
rect 186062 516218 186146 516454
rect 186382 516218 186414 516454
rect 185794 516134 186414 516218
rect 185794 515898 185826 516134
rect 186062 515898 186146 516134
rect 186382 515898 186414 516134
rect 221794 516218 221826 516454
rect 222062 516218 222146 516454
rect 222382 516218 222414 516454
rect 221794 516134 222414 516218
rect 221794 515898 221826 516134
rect 222062 515898 222146 516134
rect 222382 515898 222414 516134
rect 257794 516218 257826 516454
rect 258062 516218 258146 516454
rect 258382 516218 258414 516454
rect 257794 516134 258414 516218
rect 257794 515898 257826 516134
rect 258062 515898 258146 516134
rect 258382 515898 258414 516134
rect 293794 516218 293826 516454
rect 294062 516218 294146 516454
rect 294382 516218 294414 516454
rect 293794 516134 294414 516218
rect 293794 515898 293826 516134
rect 294062 515898 294146 516134
rect 294382 515898 294414 516134
rect 329794 516218 329826 516454
rect 330062 516218 330146 516454
rect 330382 516218 330414 516454
rect 329794 516134 330414 516218
rect 329794 515898 329826 516134
rect 330062 515898 330146 516134
rect 330382 515898 330414 516134
rect 365794 516218 365826 516454
rect 366062 516218 366146 516454
rect 366382 516218 366414 516454
rect 365794 516134 366414 516218
rect 365794 515898 365826 516134
rect 366062 515898 366146 516134
rect 366382 515898 366414 516134
rect 401794 516218 401826 516454
rect 402062 516218 402146 516454
rect 402382 516218 402414 516454
rect 401794 516134 402414 516218
rect 401794 515898 401826 516134
rect 402062 515898 402146 516134
rect 402382 515898 402414 516134
rect 570318 516218 570350 516454
rect 570586 516218 570670 516454
rect 570906 516218 570938 516454
rect 570318 516134 570938 516218
rect 570318 515898 570350 516134
rect 570586 515898 570670 516134
rect 570906 515898 570938 516134
rect -2006 480454 -1386 515898
rect 582294 484954 582914 520398
rect 23794 484718 23826 484954
rect 24062 484718 24146 484954
rect 24382 484718 24414 484954
rect 23794 484634 24414 484718
rect 23794 484398 23826 484634
rect 24062 484398 24146 484634
rect 24382 484398 24414 484634
rect 59794 484718 59826 484954
rect 60062 484718 60146 484954
rect 60382 484718 60414 484954
rect 59794 484634 60414 484718
rect 59794 484398 59826 484634
rect 60062 484398 60146 484634
rect 60382 484398 60414 484634
rect 95794 484718 95826 484954
rect 96062 484718 96146 484954
rect 96382 484718 96414 484954
rect 95794 484634 96414 484718
rect 95794 484398 95826 484634
rect 96062 484398 96146 484634
rect 96382 484398 96414 484634
rect 131794 484718 131826 484954
rect 132062 484718 132146 484954
rect 132382 484718 132414 484954
rect 131794 484634 132414 484718
rect 131794 484398 131826 484634
rect 132062 484398 132146 484634
rect 132382 484398 132414 484634
rect 167794 484718 167826 484954
rect 168062 484718 168146 484954
rect 168382 484718 168414 484954
rect 167794 484634 168414 484718
rect 167794 484398 167826 484634
rect 168062 484398 168146 484634
rect 168382 484398 168414 484634
rect 203794 484718 203826 484954
rect 204062 484718 204146 484954
rect 204382 484718 204414 484954
rect 203794 484634 204414 484718
rect 203794 484398 203826 484634
rect 204062 484398 204146 484634
rect 204382 484398 204414 484634
rect 239794 484718 239826 484954
rect 240062 484718 240146 484954
rect 240382 484718 240414 484954
rect 239794 484634 240414 484718
rect 239794 484398 239826 484634
rect 240062 484398 240146 484634
rect 240382 484398 240414 484634
rect 275794 484718 275826 484954
rect 276062 484718 276146 484954
rect 276382 484718 276414 484954
rect 275794 484634 276414 484718
rect 275794 484398 275826 484634
rect 276062 484398 276146 484634
rect 276382 484398 276414 484634
rect 311794 484718 311826 484954
rect 312062 484718 312146 484954
rect 312382 484718 312414 484954
rect 311794 484634 312414 484718
rect 311794 484398 311826 484634
rect 312062 484398 312146 484634
rect 312382 484398 312414 484634
rect 347794 484718 347826 484954
rect 348062 484718 348146 484954
rect 348382 484718 348414 484954
rect 347794 484634 348414 484718
rect 347794 484398 347826 484634
rect 348062 484398 348146 484634
rect 348382 484398 348414 484634
rect 383794 484718 383826 484954
rect 384062 484718 384146 484954
rect 384382 484718 384414 484954
rect 383794 484634 384414 484718
rect 383794 484398 383826 484634
rect 384062 484398 384146 484634
rect 384382 484398 384414 484634
rect 419794 484718 419826 484954
rect 420062 484718 420146 484954
rect 420382 484718 420414 484954
rect 419794 484634 420414 484718
rect 419794 484398 419826 484634
rect 420062 484398 420146 484634
rect 420382 484398 420414 484634
rect 455794 484718 455826 484954
rect 456062 484718 456146 484954
rect 456382 484718 456414 484954
rect 455794 484634 456414 484718
rect 455794 484398 455826 484634
rect 456062 484398 456146 484634
rect 456382 484398 456414 484634
rect 491794 484718 491826 484954
rect 492062 484718 492146 484954
rect 492382 484718 492414 484954
rect 491794 484634 492414 484718
rect 491794 484398 491826 484634
rect 492062 484398 492146 484634
rect 492382 484398 492414 484634
rect 527794 484718 527826 484954
rect 528062 484718 528146 484954
rect 528382 484718 528414 484954
rect 527794 484634 528414 484718
rect 527794 484398 527826 484634
rect 528062 484398 528146 484634
rect 528382 484398 528414 484634
rect 563794 484718 563826 484954
rect 564062 484718 564146 484954
rect 564382 484718 564414 484954
rect 563794 484634 564414 484718
rect 563794 484398 563826 484634
rect 564062 484398 564146 484634
rect 564382 484398 564414 484634
rect 582294 484718 582326 484954
rect 582562 484718 582646 484954
rect 582882 484718 582914 484954
rect 582294 484634 582914 484718
rect 582294 484398 582326 484634
rect 582562 484398 582646 484634
rect 582882 484398 582914 484634
rect -2006 480218 -1974 480454
rect -1738 480218 -1654 480454
rect -1418 480218 -1386 480454
rect -2006 480134 -1386 480218
rect -2006 479898 -1974 480134
rect -1738 479898 -1654 480134
rect -1418 479898 -1386 480134
rect 5794 480218 5826 480454
rect 6062 480218 6146 480454
rect 6382 480218 6414 480454
rect 5794 480134 6414 480218
rect 5794 479898 5826 480134
rect 6062 479898 6146 480134
rect 6382 479898 6414 480134
rect 41794 480218 41826 480454
rect 42062 480218 42146 480454
rect 42382 480218 42414 480454
rect 41794 480134 42414 480218
rect 41794 479898 41826 480134
rect 42062 479898 42146 480134
rect 42382 479898 42414 480134
rect 77794 480218 77826 480454
rect 78062 480218 78146 480454
rect 78382 480218 78414 480454
rect 77794 480134 78414 480218
rect 77794 479898 77826 480134
rect 78062 479898 78146 480134
rect 78382 479898 78414 480134
rect 113794 480218 113826 480454
rect 114062 480218 114146 480454
rect 114382 480218 114414 480454
rect 113794 480134 114414 480218
rect 113794 479898 113826 480134
rect 114062 479898 114146 480134
rect 114382 479898 114414 480134
rect 149794 480218 149826 480454
rect 150062 480218 150146 480454
rect 150382 480218 150414 480454
rect 149794 480134 150414 480218
rect 149794 479898 149826 480134
rect 150062 479898 150146 480134
rect 150382 479898 150414 480134
rect 185794 480218 185826 480454
rect 186062 480218 186146 480454
rect 186382 480218 186414 480454
rect 185794 480134 186414 480218
rect 185794 479898 185826 480134
rect 186062 479898 186146 480134
rect 186382 479898 186414 480134
rect 221794 480218 221826 480454
rect 222062 480218 222146 480454
rect 222382 480218 222414 480454
rect 221794 480134 222414 480218
rect 221794 479898 221826 480134
rect 222062 479898 222146 480134
rect 222382 479898 222414 480134
rect 257794 480218 257826 480454
rect 258062 480218 258146 480454
rect 258382 480218 258414 480454
rect 257794 480134 258414 480218
rect 257794 479898 257826 480134
rect 258062 479898 258146 480134
rect 258382 479898 258414 480134
rect 293794 480218 293826 480454
rect 294062 480218 294146 480454
rect 294382 480218 294414 480454
rect 293794 480134 294414 480218
rect 293794 479898 293826 480134
rect 294062 479898 294146 480134
rect 294382 479898 294414 480134
rect 329794 480218 329826 480454
rect 330062 480218 330146 480454
rect 330382 480218 330414 480454
rect 329794 480134 330414 480218
rect 329794 479898 329826 480134
rect 330062 479898 330146 480134
rect 330382 479898 330414 480134
rect 365794 480218 365826 480454
rect 366062 480218 366146 480454
rect 366382 480218 366414 480454
rect 365794 480134 366414 480218
rect 365794 479898 365826 480134
rect 366062 479898 366146 480134
rect 366382 479898 366414 480134
rect 401794 480218 401826 480454
rect 402062 480218 402146 480454
rect 402382 480218 402414 480454
rect 401794 480134 402414 480218
rect 401794 479898 401826 480134
rect 402062 479898 402146 480134
rect 402382 479898 402414 480134
rect 437794 480218 437826 480454
rect 438062 480218 438146 480454
rect 438382 480218 438414 480454
rect 437794 480134 438414 480218
rect 437794 479898 437826 480134
rect 438062 479898 438146 480134
rect 438382 479898 438414 480134
rect 473794 480218 473826 480454
rect 474062 480218 474146 480454
rect 474382 480218 474414 480454
rect 473794 480134 474414 480218
rect 473794 479898 473826 480134
rect 474062 479898 474146 480134
rect 474382 479898 474414 480134
rect 509794 480218 509826 480454
rect 510062 480218 510146 480454
rect 510382 480218 510414 480454
rect 509794 480134 510414 480218
rect 509794 479898 509826 480134
rect 510062 479898 510146 480134
rect 510382 479898 510414 480134
rect 545794 480218 545826 480454
rect 546062 480218 546146 480454
rect 546382 480218 546414 480454
rect 545794 480134 546414 480218
rect 545794 479898 545826 480134
rect 546062 479898 546146 480134
rect 546382 479898 546414 480134
rect -2006 444454 -1386 479898
rect 582294 448954 582914 484398
rect 13166 448718 13198 448954
rect 13434 448718 13518 448954
rect 13754 448718 13786 448954
rect 13166 448634 13786 448718
rect 13166 448398 13198 448634
rect 13434 448398 13518 448634
rect 13754 448398 13786 448634
rect 167794 448718 167826 448954
rect 168062 448718 168146 448954
rect 168382 448718 168414 448954
rect 167794 448634 168414 448718
rect 167794 448398 167826 448634
rect 168062 448398 168146 448634
rect 168382 448398 168414 448634
rect 203794 448718 203826 448954
rect 204062 448718 204146 448954
rect 204382 448718 204414 448954
rect 203794 448634 204414 448718
rect 203794 448398 203826 448634
rect 204062 448398 204146 448634
rect 204382 448398 204414 448634
rect 239794 448718 239826 448954
rect 240062 448718 240146 448954
rect 240382 448718 240414 448954
rect 239794 448634 240414 448718
rect 239794 448398 239826 448634
rect 240062 448398 240146 448634
rect 240382 448398 240414 448634
rect 275794 448718 275826 448954
rect 276062 448718 276146 448954
rect 276382 448718 276414 448954
rect 275794 448634 276414 448718
rect 275794 448398 275826 448634
rect 276062 448398 276146 448634
rect 276382 448398 276414 448634
rect 311794 448718 311826 448954
rect 312062 448718 312146 448954
rect 312382 448718 312414 448954
rect 311794 448634 312414 448718
rect 311794 448398 311826 448634
rect 312062 448398 312146 448634
rect 312382 448398 312414 448634
rect 347794 448718 347826 448954
rect 348062 448718 348146 448954
rect 348382 448718 348414 448954
rect 347794 448634 348414 448718
rect 347794 448398 347826 448634
rect 348062 448398 348146 448634
rect 348382 448398 348414 448634
rect 383794 448718 383826 448954
rect 384062 448718 384146 448954
rect 384382 448718 384414 448954
rect 383794 448634 384414 448718
rect 383794 448398 383826 448634
rect 384062 448398 384146 448634
rect 384382 448398 384414 448634
rect 419794 448718 419826 448954
rect 420062 448718 420146 448954
rect 420382 448718 420414 448954
rect 419794 448634 420414 448718
rect 419794 448398 419826 448634
rect 420062 448398 420146 448634
rect 420382 448398 420414 448634
rect 563794 448718 563826 448954
rect 564062 448718 564146 448954
rect 564382 448718 564414 448954
rect 563794 448634 564414 448718
rect 563794 448398 563826 448634
rect 564062 448398 564146 448634
rect 564382 448398 564414 448634
rect 582294 448718 582326 448954
rect 582562 448718 582646 448954
rect 582882 448718 582914 448954
rect 582294 448634 582914 448718
rect 582294 448398 582326 448634
rect 582562 448398 582646 448634
rect 582882 448398 582914 448634
rect -2006 444218 -1974 444454
rect -1738 444218 -1654 444454
rect -1418 444218 -1386 444454
rect -2006 444134 -1386 444218
rect -2006 443898 -1974 444134
rect -1738 443898 -1654 444134
rect -1418 443898 -1386 444134
rect 5794 444218 5826 444454
rect 6062 444218 6146 444454
rect 6382 444218 6414 444454
rect 5794 444134 6414 444218
rect 5794 443898 5826 444134
rect 6062 443898 6146 444134
rect 6382 443898 6414 444134
rect 185794 444218 185826 444454
rect 186062 444218 186146 444454
rect 186382 444218 186414 444454
rect 185794 444134 186414 444218
rect 185794 443898 185826 444134
rect 186062 443898 186146 444134
rect 186382 443898 186414 444134
rect 221794 444218 221826 444454
rect 222062 444218 222146 444454
rect 222382 444218 222414 444454
rect 221794 444134 222414 444218
rect 221794 443898 221826 444134
rect 222062 443898 222146 444134
rect 222382 443898 222414 444134
rect 257794 444218 257826 444454
rect 258062 444218 258146 444454
rect 258382 444218 258414 444454
rect 257794 444134 258414 444218
rect 257794 443898 257826 444134
rect 258062 443898 258146 444134
rect 258382 443898 258414 444134
rect 293794 444218 293826 444454
rect 294062 444218 294146 444454
rect 294382 444218 294414 444454
rect 293794 444134 294414 444218
rect 293794 443898 293826 444134
rect 294062 443898 294146 444134
rect 294382 443898 294414 444134
rect 329794 444218 329826 444454
rect 330062 444218 330146 444454
rect 330382 444218 330414 444454
rect 329794 444134 330414 444218
rect 329794 443898 329826 444134
rect 330062 443898 330146 444134
rect 330382 443898 330414 444134
rect 365794 444218 365826 444454
rect 366062 444218 366146 444454
rect 366382 444218 366414 444454
rect 365794 444134 366414 444218
rect 365794 443898 365826 444134
rect 366062 443898 366146 444134
rect 366382 443898 366414 444134
rect 401794 444218 401826 444454
rect 402062 444218 402146 444454
rect 402382 444218 402414 444454
rect 401794 444134 402414 444218
rect 401794 443898 401826 444134
rect 402062 443898 402146 444134
rect 402382 443898 402414 444134
rect 570318 444218 570350 444454
rect 570586 444218 570670 444454
rect 570906 444218 570938 444454
rect 570318 444134 570938 444218
rect 570318 443898 570350 444134
rect 570586 443898 570670 444134
rect 570906 443898 570938 444134
rect -2006 408454 -1386 443898
rect 582294 412954 582914 448398
rect 13166 412718 13198 412954
rect 13434 412718 13518 412954
rect 13754 412718 13786 412954
rect 13166 412634 13786 412718
rect 13166 412398 13198 412634
rect 13434 412398 13518 412634
rect 13754 412398 13786 412634
rect 167794 412718 167826 412954
rect 168062 412718 168146 412954
rect 168382 412718 168414 412954
rect 167794 412634 168414 412718
rect 167794 412398 167826 412634
rect 168062 412398 168146 412634
rect 168382 412398 168414 412634
rect 203794 412718 203826 412954
rect 204062 412718 204146 412954
rect 204382 412718 204414 412954
rect 203794 412634 204414 412718
rect 203794 412398 203826 412634
rect 204062 412398 204146 412634
rect 204382 412398 204414 412634
rect 239794 412718 239826 412954
rect 240062 412718 240146 412954
rect 240382 412718 240414 412954
rect 239794 412634 240414 412718
rect 239794 412398 239826 412634
rect 240062 412398 240146 412634
rect 240382 412398 240414 412634
rect 275794 412718 275826 412954
rect 276062 412718 276146 412954
rect 276382 412718 276414 412954
rect 275794 412634 276414 412718
rect 275794 412398 275826 412634
rect 276062 412398 276146 412634
rect 276382 412398 276414 412634
rect 311794 412718 311826 412954
rect 312062 412718 312146 412954
rect 312382 412718 312414 412954
rect 311794 412634 312414 412718
rect 311794 412398 311826 412634
rect 312062 412398 312146 412634
rect 312382 412398 312414 412634
rect 347794 412718 347826 412954
rect 348062 412718 348146 412954
rect 348382 412718 348414 412954
rect 347794 412634 348414 412718
rect 347794 412398 347826 412634
rect 348062 412398 348146 412634
rect 348382 412398 348414 412634
rect 383794 412718 383826 412954
rect 384062 412718 384146 412954
rect 384382 412718 384414 412954
rect 383794 412634 384414 412718
rect 383794 412398 383826 412634
rect 384062 412398 384146 412634
rect 384382 412398 384414 412634
rect 419794 412718 419826 412954
rect 420062 412718 420146 412954
rect 420382 412718 420414 412954
rect 419794 412634 420414 412718
rect 419794 412398 419826 412634
rect 420062 412398 420146 412634
rect 420382 412398 420414 412634
rect 563794 412718 563826 412954
rect 564062 412718 564146 412954
rect 564382 412718 564414 412954
rect 563794 412634 564414 412718
rect 563794 412398 563826 412634
rect 564062 412398 564146 412634
rect 564382 412398 564414 412634
rect 582294 412718 582326 412954
rect 582562 412718 582646 412954
rect 582882 412718 582914 412954
rect 582294 412634 582914 412718
rect 582294 412398 582326 412634
rect 582562 412398 582646 412634
rect 582882 412398 582914 412634
rect -2006 408218 -1974 408454
rect -1738 408218 -1654 408454
rect -1418 408218 -1386 408454
rect -2006 408134 -1386 408218
rect -2006 407898 -1974 408134
rect -1738 407898 -1654 408134
rect -1418 407898 -1386 408134
rect 5794 408218 5826 408454
rect 6062 408218 6146 408454
rect 6382 408218 6414 408454
rect 5794 408134 6414 408218
rect 5794 407898 5826 408134
rect 6062 407898 6146 408134
rect 6382 407898 6414 408134
rect 185794 408218 185826 408454
rect 186062 408218 186146 408454
rect 186382 408218 186414 408454
rect 185794 408134 186414 408218
rect 185794 407898 185826 408134
rect 186062 407898 186146 408134
rect 186382 407898 186414 408134
rect 221794 408218 221826 408454
rect 222062 408218 222146 408454
rect 222382 408218 222414 408454
rect 221794 408134 222414 408218
rect 221794 407898 221826 408134
rect 222062 407898 222146 408134
rect 222382 407898 222414 408134
rect 257794 408218 257826 408454
rect 258062 408218 258146 408454
rect 258382 408218 258414 408454
rect 257794 408134 258414 408218
rect 257794 407898 257826 408134
rect 258062 407898 258146 408134
rect 258382 407898 258414 408134
rect 293794 408218 293826 408454
rect 294062 408218 294146 408454
rect 294382 408218 294414 408454
rect 293794 408134 294414 408218
rect 293794 407898 293826 408134
rect 294062 407898 294146 408134
rect 294382 407898 294414 408134
rect 329794 408218 329826 408454
rect 330062 408218 330146 408454
rect 330382 408218 330414 408454
rect 329794 408134 330414 408218
rect 329794 407898 329826 408134
rect 330062 407898 330146 408134
rect 330382 407898 330414 408134
rect 365794 408218 365826 408454
rect 366062 408218 366146 408454
rect 366382 408218 366414 408454
rect 365794 408134 366414 408218
rect 365794 407898 365826 408134
rect 366062 407898 366146 408134
rect 366382 407898 366414 408134
rect 401794 408218 401826 408454
rect 402062 408218 402146 408454
rect 402382 408218 402414 408454
rect 401794 408134 402414 408218
rect 401794 407898 401826 408134
rect 402062 407898 402146 408134
rect 402382 407898 402414 408134
rect 570318 408218 570350 408454
rect 570586 408218 570670 408454
rect 570906 408218 570938 408454
rect 570318 408134 570938 408218
rect 570318 407898 570350 408134
rect 570586 407898 570670 408134
rect 570906 407898 570938 408134
rect -2006 372454 -1386 407898
rect 582294 376954 582914 412398
rect 13166 376718 13198 376954
rect 13434 376718 13518 376954
rect 13754 376718 13786 376954
rect 13166 376634 13786 376718
rect 13166 376398 13198 376634
rect 13434 376398 13518 376634
rect 13754 376398 13786 376634
rect 167794 376718 167826 376954
rect 168062 376718 168146 376954
rect 168382 376718 168414 376954
rect 167794 376634 168414 376718
rect 167794 376398 167826 376634
rect 168062 376398 168146 376634
rect 168382 376398 168414 376634
rect 203794 376718 203826 376954
rect 204062 376718 204146 376954
rect 204382 376718 204414 376954
rect 203794 376634 204414 376718
rect 203794 376398 203826 376634
rect 204062 376398 204146 376634
rect 204382 376398 204414 376634
rect 239794 376718 239826 376954
rect 240062 376718 240146 376954
rect 240382 376718 240414 376954
rect 239794 376634 240414 376718
rect 239794 376398 239826 376634
rect 240062 376398 240146 376634
rect 240382 376398 240414 376634
rect 275794 376718 275826 376954
rect 276062 376718 276146 376954
rect 276382 376718 276414 376954
rect 275794 376634 276414 376718
rect 275794 376398 275826 376634
rect 276062 376398 276146 376634
rect 276382 376398 276414 376634
rect 311794 376718 311826 376954
rect 312062 376718 312146 376954
rect 312382 376718 312414 376954
rect 311794 376634 312414 376718
rect 311794 376398 311826 376634
rect 312062 376398 312146 376634
rect 312382 376398 312414 376634
rect 347794 376718 347826 376954
rect 348062 376718 348146 376954
rect 348382 376718 348414 376954
rect 347794 376634 348414 376718
rect 347794 376398 347826 376634
rect 348062 376398 348146 376634
rect 348382 376398 348414 376634
rect 383794 376718 383826 376954
rect 384062 376718 384146 376954
rect 384382 376718 384414 376954
rect 383794 376634 384414 376718
rect 383794 376398 383826 376634
rect 384062 376398 384146 376634
rect 384382 376398 384414 376634
rect 419794 376718 419826 376954
rect 420062 376718 420146 376954
rect 420382 376718 420414 376954
rect 419794 376634 420414 376718
rect 419794 376398 419826 376634
rect 420062 376398 420146 376634
rect 420382 376398 420414 376634
rect 563794 376718 563826 376954
rect 564062 376718 564146 376954
rect 564382 376718 564414 376954
rect 563794 376634 564414 376718
rect 563794 376398 563826 376634
rect 564062 376398 564146 376634
rect 564382 376398 564414 376634
rect 582294 376718 582326 376954
rect 582562 376718 582646 376954
rect 582882 376718 582914 376954
rect 582294 376634 582914 376718
rect 582294 376398 582326 376634
rect 582562 376398 582646 376634
rect 582882 376398 582914 376634
rect -2006 372218 -1974 372454
rect -1738 372218 -1654 372454
rect -1418 372218 -1386 372454
rect -2006 372134 -1386 372218
rect -2006 371898 -1974 372134
rect -1738 371898 -1654 372134
rect -1418 371898 -1386 372134
rect 5794 372218 5826 372454
rect 6062 372218 6146 372454
rect 6382 372218 6414 372454
rect 5794 372134 6414 372218
rect 5794 371898 5826 372134
rect 6062 371898 6146 372134
rect 6382 371898 6414 372134
rect 185794 372218 185826 372454
rect 186062 372218 186146 372454
rect 186382 372218 186414 372454
rect 185794 372134 186414 372218
rect 185794 371898 185826 372134
rect 186062 371898 186146 372134
rect 186382 371898 186414 372134
rect 221794 372218 221826 372454
rect 222062 372218 222146 372454
rect 222382 372218 222414 372454
rect 221794 372134 222414 372218
rect 221794 371898 221826 372134
rect 222062 371898 222146 372134
rect 222382 371898 222414 372134
rect 257794 372218 257826 372454
rect 258062 372218 258146 372454
rect 258382 372218 258414 372454
rect 257794 372134 258414 372218
rect 257794 371898 257826 372134
rect 258062 371898 258146 372134
rect 258382 371898 258414 372134
rect 293794 372218 293826 372454
rect 294062 372218 294146 372454
rect 294382 372218 294414 372454
rect 293794 372134 294414 372218
rect 293794 371898 293826 372134
rect 294062 371898 294146 372134
rect 294382 371898 294414 372134
rect 329794 372218 329826 372454
rect 330062 372218 330146 372454
rect 330382 372218 330414 372454
rect 329794 372134 330414 372218
rect 329794 371898 329826 372134
rect 330062 371898 330146 372134
rect 330382 371898 330414 372134
rect 365794 372218 365826 372454
rect 366062 372218 366146 372454
rect 366382 372218 366414 372454
rect 365794 372134 366414 372218
rect 365794 371898 365826 372134
rect 366062 371898 366146 372134
rect 366382 371898 366414 372134
rect 401794 372218 401826 372454
rect 402062 372218 402146 372454
rect 402382 372218 402414 372454
rect 401794 372134 402414 372218
rect 401794 371898 401826 372134
rect 402062 371898 402146 372134
rect 402382 371898 402414 372134
rect 570318 372218 570350 372454
rect 570586 372218 570670 372454
rect 570906 372218 570938 372454
rect 570318 372134 570938 372218
rect 570318 371898 570350 372134
rect 570586 371898 570670 372134
rect 570906 371898 570938 372134
rect -2006 336454 -1386 371898
rect 582294 340954 582914 376398
rect 13166 340718 13198 340954
rect 13434 340718 13518 340954
rect 13754 340718 13786 340954
rect 13166 340634 13786 340718
rect 13166 340398 13198 340634
rect 13434 340398 13518 340634
rect 13754 340398 13786 340634
rect 167794 340718 167826 340954
rect 168062 340718 168146 340954
rect 168382 340718 168414 340954
rect 167794 340634 168414 340718
rect 167794 340398 167826 340634
rect 168062 340398 168146 340634
rect 168382 340398 168414 340634
rect 203794 340718 203826 340954
rect 204062 340718 204146 340954
rect 204382 340718 204414 340954
rect 203794 340634 204414 340718
rect 203794 340398 203826 340634
rect 204062 340398 204146 340634
rect 204382 340398 204414 340634
rect 239794 340718 239826 340954
rect 240062 340718 240146 340954
rect 240382 340718 240414 340954
rect 239794 340634 240414 340718
rect 239794 340398 239826 340634
rect 240062 340398 240146 340634
rect 240382 340398 240414 340634
rect 275794 340718 275826 340954
rect 276062 340718 276146 340954
rect 276382 340718 276414 340954
rect 275794 340634 276414 340718
rect 275794 340398 275826 340634
rect 276062 340398 276146 340634
rect 276382 340398 276414 340634
rect 311794 340718 311826 340954
rect 312062 340718 312146 340954
rect 312382 340718 312414 340954
rect 311794 340634 312414 340718
rect 311794 340398 311826 340634
rect 312062 340398 312146 340634
rect 312382 340398 312414 340634
rect 347794 340718 347826 340954
rect 348062 340718 348146 340954
rect 348382 340718 348414 340954
rect 347794 340634 348414 340718
rect 347794 340398 347826 340634
rect 348062 340398 348146 340634
rect 348382 340398 348414 340634
rect 383794 340718 383826 340954
rect 384062 340718 384146 340954
rect 384382 340718 384414 340954
rect 383794 340634 384414 340718
rect 383794 340398 383826 340634
rect 384062 340398 384146 340634
rect 384382 340398 384414 340634
rect 419794 340718 419826 340954
rect 420062 340718 420146 340954
rect 420382 340718 420414 340954
rect 419794 340634 420414 340718
rect 419794 340398 419826 340634
rect 420062 340398 420146 340634
rect 420382 340398 420414 340634
rect 563794 340718 563826 340954
rect 564062 340718 564146 340954
rect 564382 340718 564414 340954
rect 563794 340634 564414 340718
rect 563794 340398 563826 340634
rect 564062 340398 564146 340634
rect 564382 340398 564414 340634
rect 582294 340718 582326 340954
rect 582562 340718 582646 340954
rect 582882 340718 582914 340954
rect 582294 340634 582914 340718
rect 582294 340398 582326 340634
rect 582562 340398 582646 340634
rect 582882 340398 582914 340634
rect -2006 336218 -1974 336454
rect -1738 336218 -1654 336454
rect -1418 336218 -1386 336454
rect -2006 336134 -1386 336218
rect -2006 335898 -1974 336134
rect -1738 335898 -1654 336134
rect -1418 335898 -1386 336134
rect 5794 336218 5826 336454
rect 6062 336218 6146 336454
rect 6382 336218 6414 336454
rect 5794 336134 6414 336218
rect 5794 335898 5826 336134
rect 6062 335898 6146 336134
rect 6382 335898 6414 336134
rect 185794 336218 185826 336454
rect 186062 336218 186146 336454
rect 186382 336218 186414 336454
rect 185794 336134 186414 336218
rect 185794 335898 185826 336134
rect 186062 335898 186146 336134
rect 186382 335898 186414 336134
rect 221794 336218 221826 336454
rect 222062 336218 222146 336454
rect 222382 336218 222414 336454
rect 221794 336134 222414 336218
rect 221794 335898 221826 336134
rect 222062 335898 222146 336134
rect 222382 335898 222414 336134
rect 257794 336218 257826 336454
rect 258062 336218 258146 336454
rect 258382 336218 258414 336454
rect 257794 336134 258414 336218
rect 257794 335898 257826 336134
rect 258062 335898 258146 336134
rect 258382 335898 258414 336134
rect 293794 336218 293826 336454
rect 294062 336218 294146 336454
rect 294382 336218 294414 336454
rect 293794 336134 294414 336218
rect 293794 335898 293826 336134
rect 294062 335898 294146 336134
rect 294382 335898 294414 336134
rect 329794 336218 329826 336454
rect 330062 336218 330146 336454
rect 330382 336218 330414 336454
rect 329794 336134 330414 336218
rect 329794 335898 329826 336134
rect 330062 335898 330146 336134
rect 330382 335898 330414 336134
rect 365794 336218 365826 336454
rect 366062 336218 366146 336454
rect 366382 336218 366414 336454
rect 365794 336134 366414 336218
rect 365794 335898 365826 336134
rect 366062 335898 366146 336134
rect 366382 335898 366414 336134
rect 401794 336218 401826 336454
rect 402062 336218 402146 336454
rect 402382 336218 402414 336454
rect 401794 336134 402414 336218
rect 401794 335898 401826 336134
rect 402062 335898 402146 336134
rect 402382 335898 402414 336134
rect 570318 336218 570350 336454
rect 570586 336218 570670 336454
rect 570906 336218 570938 336454
rect 570318 336134 570938 336218
rect 570318 335898 570350 336134
rect 570586 335898 570670 336134
rect 570906 335898 570938 336134
rect -2006 300454 -1386 335898
rect 582294 304954 582914 340398
rect 13166 304718 13198 304954
rect 13434 304718 13518 304954
rect 13754 304718 13786 304954
rect 13166 304634 13786 304718
rect 13166 304398 13198 304634
rect 13434 304398 13518 304634
rect 13754 304398 13786 304634
rect 167794 304718 167826 304954
rect 168062 304718 168146 304954
rect 168382 304718 168414 304954
rect 167794 304634 168414 304718
rect 167794 304398 167826 304634
rect 168062 304398 168146 304634
rect 168382 304398 168414 304634
rect 203794 304718 203826 304954
rect 204062 304718 204146 304954
rect 204382 304718 204414 304954
rect 203794 304634 204414 304718
rect 203794 304398 203826 304634
rect 204062 304398 204146 304634
rect 204382 304398 204414 304634
rect 239794 304718 239826 304954
rect 240062 304718 240146 304954
rect 240382 304718 240414 304954
rect 239794 304634 240414 304718
rect 239794 304398 239826 304634
rect 240062 304398 240146 304634
rect 240382 304398 240414 304634
rect 275794 304718 275826 304954
rect 276062 304718 276146 304954
rect 276382 304718 276414 304954
rect 275794 304634 276414 304718
rect 275794 304398 275826 304634
rect 276062 304398 276146 304634
rect 276382 304398 276414 304634
rect 311794 304718 311826 304954
rect 312062 304718 312146 304954
rect 312382 304718 312414 304954
rect 311794 304634 312414 304718
rect 311794 304398 311826 304634
rect 312062 304398 312146 304634
rect 312382 304398 312414 304634
rect 347794 304718 347826 304954
rect 348062 304718 348146 304954
rect 348382 304718 348414 304954
rect 347794 304634 348414 304718
rect 347794 304398 347826 304634
rect 348062 304398 348146 304634
rect 348382 304398 348414 304634
rect 383794 304718 383826 304954
rect 384062 304718 384146 304954
rect 384382 304718 384414 304954
rect 383794 304634 384414 304718
rect 383794 304398 383826 304634
rect 384062 304398 384146 304634
rect 384382 304398 384414 304634
rect 419794 304718 419826 304954
rect 420062 304718 420146 304954
rect 420382 304718 420414 304954
rect 419794 304634 420414 304718
rect 419794 304398 419826 304634
rect 420062 304398 420146 304634
rect 420382 304398 420414 304634
rect 563794 304718 563826 304954
rect 564062 304718 564146 304954
rect 564382 304718 564414 304954
rect 563794 304634 564414 304718
rect 563794 304398 563826 304634
rect 564062 304398 564146 304634
rect 564382 304398 564414 304634
rect 582294 304718 582326 304954
rect 582562 304718 582646 304954
rect 582882 304718 582914 304954
rect 582294 304634 582914 304718
rect 582294 304398 582326 304634
rect 582562 304398 582646 304634
rect 582882 304398 582914 304634
rect -2006 300218 -1974 300454
rect -1738 300218 -1654 300454
rect -1418 300218 -1386 300454
rect -2006 300134 -1386 300218
rect -2006 299898 -1974 300134
rect -1738 299898 -1654 300134
rect -1418 299898 -1386 300134
rect 5794 300218 5826 300454
rect 6062 300218 6146 300454
rect 6382 300218 6414 300454
rect 5794 300134 6414 300218
rect 5794 299898 5826 300134
rect 6062 299898 6146 300134
rect 6382 299898 6414 300134
rect 185794 300218 185826 300454
rect 186062 300218 186146 300454
rect 186382 300218 186414 300454
rect 185794 300134 186414 300218
rect 185794 299898 185826 300134
rect 186062 299898 186146 300134
rect 186382 299898 186414 300134
rect 221794 300218 221826 300454
rect 222062 300218 222146 300454
rect 222382 300218 222414 300454
rect 221794 300134 222414 300218
rect 221794 299898 221826 300134
rect 222062 299898 222146 300134
rect 222382 299898 222414 300134
rect 257794 300218 257826 300454
rect 258062 300218 258146 300454
rect 258382 300218 258414 300454
rect 257794 300134 258414 300218
rect 257794 299898 257826 300134
rect 258062 299898 258146 300134
rect 258382 299898 258414 300134
rect 293794 300218 293826 300454
rect 294062 300218 294146 300454
rect 294382 300218 294414 300454
rect 293794 300134 294414 300218
rect 293794 299898 293826 300134
rect 294062 299898 294146 300134
rect 294382 299898 294414 300134
rect 329794 300218 329826 300454
rect 330062 300218 330146 300454
rect 330382 300218 330414 300454
rect 329794 300134 330414 300218
rect 329794 299898 329826 300134
rect 330062 299898 330146 300134
rect 330382 299898 330414 300134
rect 365794 300218 365826 300454
rect 366062 300218 366146 300454
rect 366382 300218 366414 300454
rect 365794 300134 366414 300218
rect 365794 299898 365826 300134
rect 366062 299898 366146 300134
rect 366382 299898 366414 300134
rect 401794 300218 401826 300454
rect 402062 300218 402146 300454
rect 402382 300218 402414 300454
rect 401794 300134 402414 300218
rect 401794 299898 401826 300134
rect 402062 299898 402146 300134
rect 402382 299898 402414 300134
rect 570318 300218 570350 300454
rect 570586 300218 570670 300454
rect 570906 300218 570938 300454
rect 570318 300134 570938 300218
rect 570318 299898 570350 300134
rect 570586 299898 570670 300134
rect 570906 299898 570938 300134
rect -2006 264454 -1386 299898
rect 582294 268954 582914 304398
rect 13166 268718 13198 268954
rect 13434 268718 13518 268954
rect 13754 268718 13786 268954
rect 13166 268634 13786 268718
rect 13166 268398 13198 268634
rect 13434 268398 13518 268634
rect 13754 268398 13786 268634
rect 167794 268718 167826 268954
rect 168062 268718 168146 268954
rect 168382 268718 168414 268954
rect 167794 268634 168414 268718
rect 167794 268398 167826 268634
rect 168062 268398 168146 268634
rect 168382 268398 168414 268634
rect 203794 268718 203826 268954
rect 204062 268718 204146 268954
rect 204382 268718 204414 268954
rect 203794 268634 204414 268718
rect 203794 268398 203826 268634
rect 204062 268398 204146 268634
rect 204382 268398 204414 268634
rect 239794 268718 239826 268954
rect 240062 268718 240146 268954
rect 240382 268718 240414 268954
rect 239794 268634 240414 268718
rect 239794 268398 239826 268634
rect 240062 268398 240146 268634
rect 240382 268398 240414 268634
rect 275794 268718 275826 268954
rect 276062 268718 276146 268954
rect 276382 268718 276414 268954
rect 275794 268634 276414 268718
rect 275794 268398 275826 268634
rect 276062 268398 276146 268634
rect 276382 268398 276414 268634
rect 311794 268718 311826 268954
rect 312062 268718 312146 268954
rect 312382 268718 312414 268954
rect 311794 268634 312414 268718
rect 311794 268398 311826 268634
rect 312062 268398 312146 268634
rect 312382 268398 312414 268634
rect 347794 268718 347826 268954
rect 348062 268718 348146 268954
rect 348382 268718 348414 268954
rect 347794 268634 348414 268718
rect 347794 268398 347826 268634
rect 348062 268398 348146 268634
rect 348382 268398 348414 268634
rect 383794 268718 383826 268954
rect 384062 268718 384146 268954
rect 384382 268718 384414 268954
rect 383794 268634 384414 268718
rect 383794 268398 383826 268634
rect 384062 268398 384146 268634
rect 384382 268398 384414 268634
rect 419794 268718 419826 268954
rect 420062 268718 420146 268954
rect 420382 268718 420414 268954
rect 419794 268634 420414 268718
rect 419794 268398 419826 268634
rect 420062 268398 420146 268634
rect 420382 268398 420414 268634
rect 563794 268718 563826 268954
rect 564062 268718 564146 268954
rect 564382 268718 564414 268954
rect 563794 268634 564414 268718
rect 563794 268398 563826 268634
rect 564062 268398 564146 268634
rect 564382 268398 564414 268634
rect 582294 268718 582326 268954
rect 582562 268718 582646 268954
rect 582882 268718 582914 268954
rect 582294 268634 582914 268718
rect 582294 268398 582326 268634
rect 582562 268398 582646 268634
rect 582882 268398 582914 268634
rect -2006 264218 -1974 264454
rect -1738 264218 -1654 264454
rect -1418 264218 -1386 264454
rect -2006 264134 -1386 264218
rect -2006 263898 -1974 264134
rect -1738 263898 -1654 264134
rect -1418 263898 -1386 264134
rect 5794 264218 5826 264454
rect 6062 264218 6146 264454
rect 6382 264218 6414 264454
rect 5794 264134 6414 264218
rect 5794 263898 5826 264134
rect 6062 263898 6146 264134
rect 6382 263898 6414 264134
rect 185794 264218 185826 264454
rect 186062 264218 186146 264454
rect 186382 264218 186414 264454
rect 185794 264134 186414 264218
rect 185794 263898 185826 264134
rect 186062 263898 186146 264134
rect 186382 263898 186414 264134
rect 221794 264218 221826 264454
rect 222062 264218 222146 264454
rect 222382 264218 222414 264454
rect 221794 264134 222414 264218
rect 221794 263898 221826 264134
rect 222062 263898 222146 264134
rect 222382 263898 222414 264134
rect 257794 264218 257826 264454
rect 258062 264218 258146 264454
rect 258382 264218 258414 264454
rect 257794 264134 258414 264218
rect 257794 263898 257826 264134
rect 258062 263898 258146 264134
rect 258382 263898 258414 264134
rect 293794 264218 293826 264454
rect 294062 264218 294146 264454
rect 294382 264218 294414 264454
rect 293794 264134 294414 264218
rect 293794 263898 293826 264134
rect 294062 263898 294146 264134
rect 294382 263898 294414 264134
rect 329794 264218 329826 264454
rect 330062 264218 330146 264454
rect 330382 264218 330414 264454
rect 329794 264134 330414 264218
rect 329794 263898 329826 264134
rect 330062 263898 330146 264134
rect 330382 263898 330414 264134
rect 365794 264218 365826 264454
rect 366062 264218 366146 264454
rect 366382 264218 366414 264454
rect 365794 264134 366414 264218
rect 365794 263898 365826 264134
rect 366062 263898 366146 264134
rect 366382 263898 366414 264134
rect 401794 264218 401826 264454
rect 402062 264218 402146 264454
rect 402382 264218 402414 264454
rect 401794 264134 402414 264218
rect 401794 263898 401826 264134
rect 402062 263898 402146 264134
rect 402382 263898 402414 264134
rect 570318 264218 570350 264454
rect 570586 264218 570670 264454
rect 570906 264218 570938 264454
rect 570318 264134 570938 264218
rect 570318 263898 570350 264134
rect 570586 263898 570670 264134
rect 570906 263898 570938 264134
rect -2006 228454 -1386 263898
rect 582294 232954 582914 268398
rect 23794 232718 23826 232954
rect 24062 232718 24146 232954
rect 24382 232718 24414 232954
rect 23794 232634 24414 232718
rect 23794 232398 23826 232634
rect 24062 232398 24146 232634
rect 24382 232398 24414 232634
rect 59794 232718 59826 232954
rect 60062 232718 60146 232954
rect 60382 232718 60414 232954
rect 59794 232634 60414 232718
rect 59794 232398 59826 232634
rect 60062 232398 60146 232634
rect 60382 232398 60414 232634
rect 95794 232718 95826 232954
rect 96062 232718 96146 232954
rect 96382 232718 96414 232954
rect 95794 232634 96414 232718
rect 95794 232398 95826 232634
rect 96062 232398 96146 232634
rect 96382 232398 96414 232634
rect 131794 232718 131826 232954
rect 132062 232718 132146 232954
rect 132382 232718 132414 232954
rect 131794 232634 132414 232718
rect 131794 232398 131826 232634
rect 132062 232398 132146 232634
rect 132382 232398 132414 232634
rect 167794 232718 167826 232954
rect 168062 232718 168146 232954
rect 168382 232718 168414 232954
rect 167794 232634 168414 232718
rect 167794 232398 167826 232634
rect 168062 232398 168146 232634
rect 168382 232398 168414 232634
rect 203794 232718 203826 232954
rect 204062 232718 204146 232954
rect 204382 232718 204414 232954
rect 203794 232634 204414 232718
rect 203794 232398 203826 232634
rect 204062 232398 204146 232634
rect 204382 232398 204414 232634
rect 239794 232718 239826 232954
rect 240062 232718 240146 232954
rect 240382 232718 240414 232954
rect 239794 232634 240414 232718
rect 239794 232398 239826 232634
rect 240062 232398 240146 232634
rect 240382 232398 240414 232634
rect 275794 232718 275826 232954
rect 276062 232718 276146 232954
rect 276382 232718 276414 232954
rect 275794 232634 276414 232718
rect 275794 232398 275826 232634
rect 276062 232398 276146 232634
rect 276382 232398 276414 232634
rect 311794 232718 311826 232954
rect 312062 232718 312146 232954
rect 312382 232718 312414 232954
rect 311794 232634 312414 232718
rect 311794 232398 311826 232634
rect 312062 232398 312146 232634
rect 312382 232398 312414 232634
rect 347794 232718 347826 232954
rect 348062 232718 348146 232954
rect 348382 232718 348414 232954
rect 347794 232634 348414 232718
rect 347794 232398 347826 232634
rect 348062 232398 348146 232634
rect 348382 232398 348414 232634
rect 383794 232718 383826 232954
rect 384062 232718 384146 232954
rect 384382 232718 384414 232954
rect 383794 232634 384414 232718
rect 383794 232398 383826 232634
rect 384062 232398 384146 232634
rect 384382 232398 384414 232634
rect 419794 232718 419826 232954
rect 420062 232718 420146 232954
rect 420382 232718 420414 232954
rect 419794 232634 420414 232718
rect 419794 232398 419826 232634
rect 420062 232398 420146 232634
rect 420382 232398 420414 232634
rect 455794 232718 455826 232954
rect 456062 232718 456146 232954
rect 456382 232718 456414 232954
rect 455794 232634 456414 232718
rect 455794 232398 455826 232634
rect 456062 232398 456146 232634
rect 456382 232398 456414 232634
rect 491794 232718 491826 232954
rect 492062 232718 492146 232954
rect 492382 232718 492414 232954
rect 491794 232634 492414 232718
rect 491794 232398 491826 232634
rect 492062 232398 492146 232634
rect 492382 232398 492414 232634
rect 527794 232718 527826 232954
rect 528062 232718 528146 232954
rect 528382 232718 528414 232954
rect 527794 232634 528414 232718
rect 527794 232398 527826 232634
rect 528062 232398 528146 232634
rect 528382 232398 528414 232634
rect 563794 232718 563826 232954
rect 564062 232718 564146 232954
rect 564382 232718 564414 232954
rect 563794 232634 564414 232718
rect 563794 232398 563826 232634
rect 564062 232398 564146 232634
rect 564382 232398 564414 232634
rect 582294 232718 582326 232954
rect 582562 232718 582646 232954
rect 582882 232718 582914 232954
rect 582294 232634 582914 232718
rect 582294 232398 582326 232634
rect 582562 232398 582646 232634
rect 582882 232398 582914 232634
rect -2006 228218 -1974 228454
rect -1738 228218 -1654 228454
rect -1418 228218 -1386 228454
rect -2006 228134 -1386 228218
rect -2006 227898 -1974 228134
rect -1738 227898 -1654 228134
rect -1418 227898 -1386 228134
rect 5794 228218 5826 228454
rect 6062 228218 6146 228454
rect 6382 228218 6414 228454
rect 5794 228134 6414 228218
rect 5794 227898 5826 228134
rect 6062 227898 6146 228134
rect 6382 227898 6414 228134
rect 41794 228218 41826 228454
rect 42062 228218 42146 228454
rect 42382 228218 42414 228454
rect 41794 228134 42414 228218
rect 41794 227898 41826 228134
rect 42062 227898 42146 228134
rect 42382 227898 42414 228134
rect 77794 228218 77826 228454
rect 78062 228218 78146 228454
rect 78382 228218 78414 228454
rect 77794 228134 78414 228218
rect 77794 227898 77826 228134
rect 78062 227898 78146 228134
rect 78382 227898 78414 228134
rect 113794 228218 113826 228454
rect 114062 228218 114146 228454
rect 114382 228218 114414 228454
rect 113794 228134 114414 228218
rect 113794 227898 113826 228134
rect 114062 227898 114146 228134
rect 114382 227898 114414 228134
rect 149794 228218 149826 228454
rect 150062 228218 150146 228454
rect 150382 228218 150414 228454
rect 149794 228134 150414 228218
rect 149794 227898 149826 228134
rect 150062 227898 150146 228134
rect 150382 227898 150414 228134
rect 185794 228218 185826 228454
rect 186062 228218 186146 228454
rect 186382 228218 186414 228454
rect 185794 228134 186414 228218
rect 185794 227898 185826 228134
rect 186062 227898 186146 228134
rect 186382 227898 186414 228134
rect 221794 228218 221826 228454
rect 222062 228218 222146 228454
rect 222382 228218 222414 228454
rect 221794 228134 222414 228218
rect 221794 227898 221826 228134
rect 222062 227898 222146 228134
rect 222382 227898 222414 228134
rect 257794 228218 257826 228454
rect 258062 228218 258146 228454
rect 258382 228218 258414 228454
rect 257794 228134 258414 228218
rect 257794 227898 257826 228134
rect 258062 227898 258146 228134
rect 258382 227898 258414 228134
rect 293794 228218 293826 228454
rect 294062 228218 294146 228454
rect 294382 228218 294414 228454
rect 293794 228134 294414 228218
rect 293794 227898 293826 228134
rect 294062 227898 294146 228134
rect 294382 227898 294414 228134
rect 329794 228218 329826 228454
rect 330062 228218 330146 228454
rect 330382 228218 330414 228454
rect 329794 228134 330414 228218
rect 329794 227898 329826 228134
rect 330062 227898 330146 228134
rect 330382 227898 330414 228134
rect 365794 228218 365826 228454
rect 366062 228218 366146 228454
rect 366382 228218 366414 228454
rect 365794 228134 366414 228218
rect 365794 227898 365826 228134
rect 366062 227898 366146 228134
rect 366382 227898 366414 228134
rect 401794 228218 401826 228454
rect 402062 228218 402146 228454
rect 402382 228218 402414 228454
rect 401794 228134 402414 228218
rect 401794 227898 401826 228134
rect 402062 227898 402146 228134
rect 402382 227898 402414 228134
rect 437794 228218 437826 228454
rect 438062 228218 438146 228454
rect 438382 228218 438414 228454
rect 437794 228134 438414 228218
rect 437794 227898 437826 228134
rect 438062 227898 438146 228134
rect 438382 227898 438414 228134
rect 473794 228218 473826 228454
rect 474062 228218 474146 228454
rect 474382 228218 474414 228454
rect 473794 228134 474414 228218
rect 473794 227898 473826 228134
rect 474062 227898 474146 228134
rect 474382 227898 474414 228134
rect 509794 228218 509826 228454
rect 510062 228218 510146 228454
rect 510382 228218 510414 228454
rect 509794 228134 510414 228218
rect 509794 227898 509826 228134
rect 510062 227898 510146 228134
rect 510382 227898 510414 228134
rect 545794 228218 545826 228454
rect 546062 228218 546146 228454
rect 546382 228218 546414 228454
rect 545794 228134 546414 228218
rect 545794 227898 545826 228134
rect 546062 227898 546146 228134
rect 546382 227898 546414 228134
rect -2006 192454 -1386 227898
rect 582294 196954 582914 232398
rect 13166 196718 13198 196954
rect 13434 196718 13518 196954
rect 13754 196718 13786 196954
rect 13166 196634 13786 196718
rect 13166 196398 13198 196634
rect 13434 196398 13518 196634
rect 13754 196398 13786 196634
rect 167794 196718 167826 196954
rect 168062 196718 168146 196954
rect 168382 196718 168414 196954
rect 167794 196634 168414 196718
rect 167794 196398 167826 196634
rect 168062 196398 168146 196634
rect 168382 196398 168414 196634
rect 203794 196718 203826 196954
rect 204062 196718 204146 196954
rect 204382 196718 204414 196954
rect 203794 196634 204414 196718
rect 203794 196398 203826 196634
rect 204062 196398 204146 196634
rect 204382 196398 204414 196634
rect 239794 196718 239826 196954
rect 240062 196718 240146 196954
rect 240382 196718 240414 196954
rect 239794 196634 240414 196718
rect 239794 196398 239826 196634
rect 240062 196398 240146 196634
rect 240382 196398 240414 196634
rect 275794 196718 275826 196954
rect 276062 196718 276146 196954
rect 276382 196718 276414 196954
rect 275794 196634 276414 196718
rect 275794 196398 275826 196634
rect 276062 196398 276146 196634
rect 276382 196398 276414 196634
rect 311794 196718 311826 196954
rect 312062 196718 312146 196954
rect 312382 196718 312414 196954
rect 311794 196634 312414 196718
rect 311794 196398 311826 196634
rect 312062 196398 312146 196634
rect 312382 196398 312414 196634
rect 347794 196718 347826 196954
rect 348062 196718 348146 196954
rect 348382 196718 348414 196954
rect 347794 196634 348414 196718
rect 347794 196398 347826 196634
rect 348062 196398 348146 196634
rect 348382 196398 348414 196634
rect 383794 196718 383826 196954
rect 384062 196718 384146 196954
rect 384382 196718 384414 196954
rect 383794 196634 384414 196718
rect 383794 196398 383826 196634
rect 384062 196398 384146 196634
rect 384382 196398 384414 196634
rect 419794 196718 419826 196954
rect 420062 196718 420146 196954
rect 420382 196718 420414 196954
rect 419794 196634 420414 196718
rect 419794 196398 419826 196634
rect 420062 196398 420146 196634
rect 420382 196398 420414 196634
rect 563794 196718 563826 196954
rect 564062 196718 564146 196954
rect 564382 196718 564414 196954
rect 563794 196634 564414 196718
rect 563794 196398 563826 196634
rect 564062 196398 564146 196634
rect 564382 196398 564414 196634
rect 582294 196718 582326 196954
rect 582562 196718 582646 196954
rect 582882 196718 582914 196954
rect 582294 196634 582914 196718
rect 582294 196398 582326 196634
rect 582562 196398 582646 196634
rect 582882 196398 582914 196634
rect -2006 192218 -1974 192454
rect -1738 192218 -1654 192454
rect -1418 192218 -1386 192454
rect -2006 192134 -1386 192218
rect -2006 191898 -1974 192134
rect -1738 191898 -1654 192134
rect -1418 191898 -1386 192134
rect 5794 192218 5826 192454
rect 6062 192218 6146 192454
rect 6382 192218 6414 192454
rect 5794 192134 6414 192218
rect 5794 191898 5826 192134
rect 6062 191898 6146 192134
rect 6382 191898 6414 192134
rect 185794 192218 185826 192454
rect 186062 192218 186146 192454
rect 186382 192218 186414 192454
rect 185794 192134 186414 192218
rect 185794 191898 185826 192134
rect 186062 191898 186146 192134
rect 186382 191898 186414 192134
rect 221794 192218 221826 192454
rect 222062 192218 222146 192454
rect 222382 192218 222414 192454
rect 221794 192134 222414 192218
rect 221794 191898 221826 192134
rect 222062 191898 222146 192134
rect 222382 191898 222414 192134
rect 257794 192218 257826 192454
rect 258062 192218 258146 192454
rect 258382 192218 258414 192454
rect 257794 192134 258414 192218
rect 257794 191898 257826 192134
rect 258062 191898 258146 192134
rect 258382 191898 258414 192134
rect 293794 192218 293826 192454
rect 294062 192218 294146 192454
rect 294382 192218 294414 192454
rect 293794 192134 294414 192218
rect 293794 191898 293826 192134
rect 294062 191898 294146 192134
rect 294382 191898 294414 192134
rect 329794 192218 329826 192454
rect 330062 192218 330146 192454
rect 330382 192218 330414 192454
rect 329794 192134 330414 192218
rect 329794 191898 329826 192134
rect 330062 191898 330146 192134
rect 330382 191898 330414 192134
rect 365794 192218 365826 192454
rect 366062 192218 366146 192454
rect 366382 192218 366414 192454
rect 365794 192134 366414 192218
rect 365794 191898 365826 192134
rect 366062 191898 366146 192134
rect 366382 191898 366414 192134
rect 401794 192218 401826 192454
rect 402062 192218 402146 192454
rect 402382 192218 402414 192454
rect 401794 192134 402414 192218
rect 401794 191898 401826 192134
rect 402062 191898 402146 192134
rect 402382 191898 402414 192134
rect 570318 192218 570350 192454
rect 570586 192218 570670 192454
rect 570906 192218 570938 192454
rect 570318 192134 570938 192218
rect 570318 191898 570350 192134
rect 570586 191898 570670 192134
rect 570906 191898 570938 192134
rect -2006 156454 -1386 191898
rect 582294 160954 582914 196398
rect 13166 160718 13198 160954
rect 13434 160718 13518 160954
rect 13754 160718 13786 160954
rect 13166 160634 13786 160718
rect 13166 160398 13198 160634
rect 13434 160398 13518 160634
rect 13754 160398 13786 160634
rect 167794 160718 167826 160954
rect 168062 160718 168146 160954
rect 168382 160718 168414 160954
rect 167794 160634 168414 160718
rect 167794 160398 167826 160634
rect 168062 160398 168146 160634
rect 168382 160398 168414 160634
rect 203794 160718 203826 160954
rect 204062 160718 204146 160954
rect 204382 160718 204414 160954
rect 203794 160634 204414 160718
rect 203794 160398 203826 160634
rect 204062 160398 204146 160634
rect 204382 160398 204414 160634
rect 239794 160718 239826 160954
rect 240062 160718 240146 160954
rect 240382 160718 240414 160954
rect 239794 160634 240414 160718
rect 239794 160398 239826 160634
rect 240062 160398 240146 160634
rect 240382 160398 240414 160634
rect 275794 160718 275826 160954
rect 276062 160718 276146 160954
rect 276382 160718 276414 160954
rect 275794 160634 276414 160718
rect 275794 160398 275826 160634
rect 276062 160398 276146 160634
rect 276382 160398 276414 160634
rect 311794 160718 311826 160954
rect 312062 160718 312146 160954
rect 312382 160718 312414 160954
rect 311794 160634 312414 160718
rect 311794 160398 311826 160634
rect 312062 160398 312146 160634
rect 312382 160398 312414 160634
rect 347794 160718 347826 160954
rect 348062 160718 348146 160954
rect 348382 160718 348414 160954
rect 347794 160634 348414 160718
rect 347794 160398 347826 160634
rect 348062 160398 348146 160634
rect 348382 160398 348414 160634
rect 383794 160718 383826 160954
rect 384062 160718 384146 160954
rect 384382 160718 384414 160954
rect 383794 160634 384414 160718
rect 383794 160398 383826 160634
rect 384062 160398 384146 160634
rect 384382 160398 384414 160634
rect 419794 160718 419826 160954
rect 420062 160718 420146 160954
rect 420382 160718 420414 160954
rect 419794 160634 420414 160718
rect 419794 160398 419826 160634
rect 420062 160398 420146 160634
rect 420382 160398 420414 160634
rect 563794 160718 563826 160954
rect 564062 160718 564146 160954
rect 564382 160718 564414 160954
rect 563794 160634 564414 160718
rect 563794 160398 563826 160634
rect 564062 160398 564146 160634
rect 564382 160398 564414 160634
rect 582294 160718 582326 160954
rect 582562 160718 582646 160954
rect 582882 160718 582914 160954
rect 582294 160634 582914 160718
rect 582294 160398 582326 160634
rect 582562 160398 582646 160634
rect 582882 160398 582914 160634
rect -2006 156218 -1974 156454
rect -1738 156218 -1654 156454
rect -1418 156218 -1386 156454
rect -2006 156134 -1386 156218
rect -2006 155898 -1974 156134
rect -1738 155898 -1654 156134
rect -1418 155898 -1386 156134
rect 5794 156218 5826 156454
rect 6062 156218 6146 156454
rect 6382 156218 6414 156454
rect 5794 156134 6414 156218
rect 5794 155898 5826 156134
rect 6062 155898 6146 156134
rect 6382 155898 6414 156134
rect 185794 156218 185826 156454
rect 186062 156218 186146 156454
rect 186382 156218 186414 156454
rect 185794 156134 186414 156218
rect 185794 155898 185826 156134
rect 186062 155898 186146 156134
rect 186382 155898 186414 156134
rect 221794 156218 221826 156454
rect 222062 156218 222146 156454
rect 222382 156218 222414 156454
rect 221794 156134 222414 156218
rect 221794 155898 221826 156134
rect 222062 155898 222146 156134
rect 222382 155898 222414 156134
rect 257794 156218 257826 156454
rect 258062 156218 258146 156454
rect 258382 156218 258414 156454
rect 257794 156134 258414 156218
rect 257794 155898 257826 156134
rect 258062 155898 258146 156134
rect 258382 155898 258414 156134
rect 293794 156218 293826 156454
rect 294062 156218 294146 156454
rect 294382 156218 294414 156454
rect 293794 156134 294414 156218
rect 293794 155898 293826 156134
rect 294062 155898 294146 156134
rect 294382 155898 294414 156134
rect 329794 156218 329826 156454
rect 330062 156218 330146 156454
rect 330382 156218 330414 156454
rect 329794 156134 330414 156218
rect 329794 155898 329826 156134
rect 330062 155898 330146 156134
rect 330382 155898 330414 156134
rect 365794 156218 365826 156454
rect 366062 156218 366146 156454
rect 366382 156218 366414 156454
rect 365794 156134 366414 156218
rect 365794 155898 365826 156134
rect 366062 155898 366146 156134
rect 366382 155898 366414 156134
rect 401794 156218 401826 156454
rect 402062 156218 402146 156454
rect 402382 156218 402414 156454
rect 401794 156134 402414 156218
rect 401794 155898 401826 156134
rect 402062 155898 402146 156134
rect 402382 155898 402414 156134
rect 570318 156218 570350 156454
rect 570586 156218 570670 156454
rect 570906 156218 570938 156454
rect 570318 156134 570938 156218
rect 570318 155898 570350 156134
rect 570586 155898 570670 156134
rect 570906 155898 570938 156134
rect -2006 120454 -1386 155898
rect 582294 124954 582914 160398
rect 23794 124718 23826 124954
rect 24062 124718 24146 124954
rect 24382 124718 24414 124954
rect 23794 124634 24414 124718
rect 23794 124398 23826 124634
rect 24062 124398 24146 124634
rect 24382 124398 24414 124634
rect 59794 124718 59826 124954
rect 60062 124718 60146 124954
rect 60382 124718 60414 124954
rect 59794 124634 60414 124718
rect 59794 124398 59826 124634
rect 60062 124398 60146 124634
rect 60382 124398 60414 124634
rect 95794 124718 95826 124954
rect 96062 124718 96146 124954
rect 96382 124718 96414 124954
rect 95794 124634 96414 124718
rect 95794 124398 95826 124634
rect 96062 124398 96146 124634
rect 96382 124398 96414 124634
rect 131794 124718 131826 124954
rect 132062 124718 132146 124954
rect 132382 124718 132414 124954
rect 131794 124634 132414 124718
rect 131794 124398 131826 124634
rect 132062 124398 132146 124634
rect 132382 124398 132414 124634
rect 167794 124718 167826 124954
rect 168062 124718 168146 124954
rect 168382 124718 168414 124954
rect 167794 124634 168414 124718
rect 167794 124398 167826 124634
rect 168062 124398 168146 124634
rect 168382 124398 168414 124634
rect 203794 124718 203826 124954
rect 204062 124718 204146 124954
rect 204382 124718 204414 124954
rect 203794 124634 204414 124718
rect 203794 124398 203826 124634
rect 204062 124398 204146 124634
rect 204382 124398 204414 124634
rect 239794 124718 239826 124954
rect 240062 124718 240146 124954
rect 240382 124718 240414 124954
rect 239794 124634 240414 124718
rect 239794 124398 239826 124634
rect 240062 124398 240146 124634
rect 240382 124398 240414 124634
rect 275794 124718 275826 124954
rect 276062 124718 276146 124954
rect 276382 124718 276414 124954
rect 275794 124634 276414 124718
rect 275794 124398 275826 124634
rect 276062 124398 276146 124634
rect 276382 124398 276414 124634
rect 311794 124718 311826 124954
rect 312062 124718 312146 124954
rect 312382 124718 312414 124954
rect 311794 124634 312414 124718
rect 311794 124398 311826 124634
rect 312062 124398 312146 124634
rect 312382 124398 312414 124634
rect 347794 124718 347826 124954
rect 348062 124718 348146 124954
rect 348382 124718 348414 124954
rect 347794 124634 348414 124718
rect 347794 124398 347826 124634
rect 348062 124398 348146 124634
rect 348382 124398 348414 124634
rect 383794 124718 383826 124954
rect 384062 124718 384146 124954
rect 384382 124718 384414 124954
rect 383794 124634 384414 124718
rect 383794 124398 383826 124634
rect 384062 124398 384146 124634
rect 384382 124398 384414 124634
rect 419794 124718 419826 124954
rect 420062 124718 420146 124954
rect 420382 124718 420414 124954
rect 419794 124634 420414 124718
rect 419794 124398 419826 124634
rect 420062 124398 420146 124634
rect 420382 124398 420414 124634
rect 455794 124718 455826 124954
rect 456062 124718 456146 124954
rect 456382 124718 456414 124954
rect 455794 124634 456414 124718
rect 455794 124398 455826 124634
rect 456062 124398 456146 124634
rect 456382 124398 456414 124634
rect 491794 124718 491826 124954
rect 492062 124718 492146 124954
rect 492382 124718 492414 124954
rect 491794 124634 492414 124718
rect 491794 124398 491826 124634
rect 492062 124398 492146 124634
rect 492382 124398 492414 124634
rect 527794 124718 527826 124954
rect 528062 124718 528146 124954
rect 528382 124718 528414 124954
rect 527794 124634 528414 124718
rect 527794 124398 527826 124634
rect 528062 124398 528146 124634
rect 528382 124398 528414 124634
rect 563794 124718 563826 124954
rect 564062 124718 564146 124954
rect 564382 124718 564414 124954
rect 563794 124634 564414 124718
rect 563794 124398 563826 124634
rect 564062 124398 564146 124634
rect 564382 124398 564414 124634
rect 582294 124718 582326 124954
rect 582562 124718 582646 124954
rect 582882 124718 582914 124954
rect 582294 124634 582914 124718
rect 582294 124398 582326 124634
rect 582562 124398 582646 124634
rect 582882 124398 582914 124634
rect -2006 120218 -1974 120454
rect -1738 120218 -1654 120454
rect -1418 120218 -1386 120454
rect -2006 120134 -1386 120218
rect -2006 119898 -1974 120134
rect -1738 119898 -1654 120134
rect -1418 119898 -1386 120134
rect 5794 120218 5826 120454
rect 6062 120218 6146 120454
rect 6382 120218 6414 120454
rect 5794 120134 6414 120218
rect 5794 119898 5826 120134
rect 6062 119898 6146 120134
rect 6382 119898 6414 120134
rect 41794 120218 41826 120454
rect 42062 120218 42146 120454
rect 42382 120218 42414 120454
rect 41794 120134 42414 120218
rect 41794 119898 41826 120134
rect 42062 119898 42146 120134
rect 42382 119898 42414 120134
rect 77794 120218 77826 120454
rect 78062 120218 78146 120454
rect 78382 120218 78414 120454
rect 77794 120134 78414 120218
rect 77794 119898 77826 120134
rect 78062 119898 78146 120134
rect 78382 119898 78414 120134
rect 113794 120218 113826 120454
rect 114062 120218 114146 120454
rect 114382 120218 114414 120454
rect 113794 120134 114414 120218
rect 113794 119898 113826 120134
rect 114062 119898 114146 120134
rect 114382 119898 114414 120134
rect 149794 120218 149826 120454
rect 150062 120218 150146 120454
rect 150382 120218 150414 120454
rect 149794 120134 150414 120218
rect 149794 119898 149826 120134
rect 150062 119898 150146 120134
rect 150382 119898 150414 120134
rect 185794 120218 185826 120454
rect 186062 120218 186146 120454
rect 186382 120218 186414 120454
rect 185794 120134 186414 120218
rect 185794 119898 185826 120134
rect 186062 119898 186146 120134
rect 186382 119898 186414 120134
rect 221794 120218 221826 120454
rect 222062 120218 222146 120454
rect 222382 120218 222414 120454
rect 221794 120134 222414 120218
rect 221794 119898 221826 120134
rect 222062 119898 222146 120134
rect 222382 119898 222414 120134
rect 257794 120218 257826 120454
rect 258062 120218 258146 120454
rect 258382 120218 258414 120454
rect 257794 120134 258414 120218
rect 257794 119898 257826 120134
rect 258062 119898 258146 120134
rect 258382 119898 258414 120134
rect 293794 120218 293826 120454
rect 294062 120218 294146 120454
rect 294382 120218 294414 120454
rect 293794 120134 294414 120218
rect 293794 119898 293826 120134
rect 294062 119898 294146 120134
rect 294382 119898 294414 120134
rect 329794 120218 329826 120454
rect 330062 120218 330146 120454
rect 330382 120218 330414 120454
rect 329794 120134 330414 120218
rect 329794 119898 329826 120134
rect 330062 119898 330146 120134
rect 330382 119898 330414 120134
rect 365794 120218 365826 120454
rect 366062 120218 366146 120454
rect 366382 120218 366414 120454
rect 365794 120134 366414 120218
rect 365794 119898 365826 120134
rect 366062 119898 366146 120134
rect 366382 119898 366414 120134
rect 401794 120218 401826 120454
rect 402062 120218 402146 120454
rect 402382 120218 402414 120454
rect 401794 120134 402414 120218
rect 401794 119898 401826 120134
rect 402062 119898 402146 120134
rect 402382 119898 402414 120134
rect 437794 120218 437826 120454
rect 438062 120218 438146 120454
rect 438382 120218 438414 120454
rect 437794 120134 438414 120218
rect 437794 119898 437826 120134
rect 438062 119898 438146 120134
rect 438382 119898 438414 120134
rect 473794 120218 473826 120454
rect 474062 120218 474146 120454
rect 474382 120218 474414 120454
rect 473794 120134 474414 120218
rect 473794 119898 473826 120134
rect 474062 119898 474146 120134
rect 474382 119898 474414 120134
rect 509794 120218 509826 120454
rect 510062 120218 510146 120454
rect 510382 120218 510414 120454
rect 509794 120134 510414 120218
rect 509794 119898 509826 120134
rect 510062 119898 510146 120134
rect 510382 119898 510414 120134
rect 545794 120218 545826 120454
rect 546062 120218 546146 120454
rect 546382 120218 546414 120454
rect 545794 120134 546414 120218
rect 545794 119898 545826 120134
rect 546062 119898 546146 120134
rect 546382 119898 546414 120134
rect -2006 84454 -1386 119898
rect 582294 88954 582914 124398
rect 13166 88718 13198 88954
rect 13434 88718 13518 88954
rect 13754 88718 13786 88954
rect 13166 88634 13786 88718
rect 13166 88398 13198 88634
rect 13434 88398 13518 88634
rect 13754 88398 13786 88634
rect 167794 88718 167826 88954
rect 168062 88718 168146 88954
rect 168382 88718 168414 88954
rect 167794 88634 168414 88718
rect 167794 88398 167826 88634
rect 168062 88398 168146 88634
rect 168382 88398 168414 88634
rect 291558 88718 291590 88954
rect 291826 88718 291910 88954
rect 292146 88718 292178 88954
rect 291558 88634 292178 88718
rect 291558 88398 291590 88634
rect 291826 88398 291910 88634
rect 292146 88398 292178 88634
rect 419794 88718 419826 88954
rect 420062 88718 420146 88954
rect 420382 88718 420414 88954
rect 419794 88634 420414 88718
rect 419794 88398 419826 88634
rect 420062 88398 420146 88634
rect 420382 88398 420414 88634
rect 563794 88718 563826 88954
rect 564062 88718 564146 88954
rect 564382 88718 564414 88954
rect 563794 88634 564414 88718
rect 563794 88398 563826 88634
rect 564062 88398 564146 88634
rect 564382 88398 564414 88634
rect 582294 88718 582326 88954
rect 582562 88718 582646 88954
rect 582882 88718 582914 88954
rect 582294 88634 582914 88718
rect 582294 88398 582326 88634
rect 582562 88398 582646 88634
rect 582882 88398 582914 88634
rect -2006 84218 -1974 84454
rect -1738 84218 -1654 84454
rect -1418 84218 -1386 84454
rect -2006 84134 -1386 84218
rect -2006 83898 -1974 84134
rect -1738 83898 -1654 84134
rect -1418 83898 -1386 84134
rect 5794 84218 5826 84454
rect 6062 84218 6146 84454
rect 6382 84218 6414 84454
rect 5794 84134 6414 84218
rect 5794 83898 5826 84134
rect 6062 83898 6146 84134
rect 6382 83898 6414 84134
rect 173062 84218 173094 84454
rect 173330 84218 173414 84454
rect 173650 84218 173682 84454
rect 173062 84134 173682 84218
rect 173062 83898 173094 84134
rect 173330 83898 173414 84134
rect 173650 83898 173682 84134
rect 293794 84218 293826 84454
rect 294062 84218 294146 84454
rect 294382 84218 294414 84454
rect 293794 84134 294414 84218
rect 293794 83898 293826 84134
rect 294062 83898 294146 84134
rect 294382 83898 294414 84134
rect 401794 84218 401826 84454
rect 402062 84218 402146 84454
rect 402382 84218 402414 84454
rect 401794 84134 402414 84218
rect 401794 83898 401826 84134
rect 402062 83898 402146 84134
rect 402382 83898 402414 84134
rect 570318 84218 570350 84454
rect 570586 84218 570670 84454
rect 570906 84218 570938 84454
rect 570318 84134 570938 84218
rect 570318 83898 570350 84134
rect 570586 83898 570670 84134
rect 570906 83898 570938 84134
rect -2006 48454 -1386 83898
rect 582294 52954 582914 88398
rect 13166 52718 13198 52954
rect 13434 52718 13518 52954
rect 13754 52718 13786 52954
rect 13166 52634 13786 52718
rect 13166 52398 13198 52634
rect 13434 52398 13518 52634
rect 13754 52398 13786 52634
rect 167794 52718 167826 52954
rect 168062 52718 168146 52954
rect 168382 52718 168414 52954
rect 167794 52634 168414 52718
rect 167794 52398 167826 52634
rect 168062 52398 168146 52634
rect 168382 52398 168414 52634
rect 291558 52718 291590 52954
rect 291826 52718 291910 52954
rect 292146 52718 292178 52954
rect 291558 52634 292178 52718
rect 291558 52398 291590 52634
rect 291826 52398 291910 52634
rect 292146 52398 292178 52634
rect 419794 52718 419826 52954
rect 420062 52718 420146 52954
rect 420382 52718 420414 52954
rect 419794 52634 420414 52718
rect 419794 52398 419826 52634
rect 420062 52398 420146 52634
rect 420382 52398 420414 52634
rect 563794 52718 563826 52954
rect 564062 52718 564146 52954
rect 564382 52718 564414 52954
rect 563794 52634 564414 52718
rect 563794 52398 563826 52634
rect 564062 52398 564146 52634
rect 564382 52398 564414 52634
rect 582294 52718 582326 52954
rect 582562 52718 582646 52954
rect 582882 52718 582914 52954
rect 582294 52634 582914 52718
rect 582294 52398 582326 52634
rect 582562 52398 582646 52634
rect 582882 52398 582914 52634
rect -2006 48218 -1974 48454
rect -1738 48218 -1654 48454
rect -1418 48218 -1386 48454
rect -2006 48134 -1386 48218
rect -2006 47898 -1974 48134
rect -1738 47898 -1654 48134
rect -1418 47898 -1386 48134
rect 5794 48218 5826 48454
rect 6062 48218 6146 48454
rect 6382 48218 6414 48454
rect 5794 48134 6414 48218
rect 5794 47898 5826 48134
rect 6062 47898 6146 48134
rect 6382 47898 6414 48134
rect 173062 48218 173094 48454
rect 173330 48218 173414 48454
rect 173650 48218 173682 48454
rect 173062 48134 173682 48218
rect 173062 47898 173094 48134
rect 173330 47898 173414 48134
rect 173650 47898 173682 48134
rect 293794 48218 293826 48454
rect 294062 48218 294146 48454
rect 294382 48218 294414 48454
rect 293794 48134 294414 48218
rect 293794 47898 293826 48134
rect 294062 47898 294146 48134
rect 294382 47898 294414 48134
rect 401794 48218 401826 48454
rect 402062 48218 402146 48454
rect 402382 48218 402414 48454
rect 401794 48134 402414 48218
rect 401794 47898 401826 48134
rect 402062 47898 402146 48134
rect 402382 47898 402414 48134
rect 570318 48218 570350 48454
rect 570586 48218 570670 48454
rect 570906 48218 570938 48454
rect 570318 48134 570938 48218
rect 570318 47898 570350 48134
rect 570586 47898 570670 48134
rect 570906 47898 570938 48134
rect -2006 12454 -1386 47898
rect 582294 16954 582914 52398
rect 23794 16718 23826 16954
rect 24062 16718 24146 16954
rect 24382 16718 24414 16954
rect 23794 16634 24414 16718
rect 23794 16398 23826 16634
rect 24062 16398 24146 16634
rect 24382 16398 24414 16634
rect 59794 16718 59826 16954
rect 60062 16718 60146 16954
rect 60382 16718 60414 16954
rect 59794 16634 60414 16718
rect 59794 16398 59826 16634
rect 60062 16398 60146 16634
rect 60382 16398 60414 16634
rect 95794 16718 95826 16954
rect 96062 16718 96146 16954
rect 96382 16718 96414 16954
rect 95794 16634 96414 16718
rect 95794 16398 95826 16634
rect 96062 16398 96146 16634
rect 96382 16398 96414 16634
rect 131794 16718 131826 16954
rect 132062 16718 132146 16954
rect 132382 16718 132414 16954
rect 131794 16634 132414 16718
rect 131794 16398 131826 16634
rect 132062 16398 132146 16634
rect 132382 16398 132414 16634
rect 167794 16718 167826 16954
rect 168062 16718 168146 16954
rect 168382 16718 168414 16954
rect 167794 16634 168414 16718
rect 167794 16398 167826 16634
rect 168062 16398 168146 16634
rect 168382 16398 168414 16634
rect 203794 16718 203826 16954
rect 204062 16718 204146 16954
rect 204382 16718 204414 16954
rect 203794 16634 204414 16718
rect 203794 16398 203826 16634
rect 204062 16398 204146 16634
rect 204382 16398 204414 16634
rect 239794 16718 239826 16954
rect 240062 16718 240146 16954
rect 240382 16718 240414 16954
rect 239794 16634 240414 16718
rect 239794 16398 239826 16634
rect 240062 16398 240146 16634
rect 240382 16398 240414 16634
rect 275794 16718 275826 16954
rect 276062 16718 276146 16954
rect 276382 16718 276414 16954
rect 275794 16634 276414 16718
rect 275794 16398 275826 16634
rect 276062 16398 276146 16634
rect 276382 16398 276414 16634
rect 311794 16718 311826 16954
rect 312062 16718 312146 16954
rect 312382 16718 312414 16954
rect 311794 16634 312414 16718
rect 311794 16398 311826 16634
rect 312062 16398 312146 16634
rect 312382 16398 312414 16634
rect 347794 16718 347826 16954
rect 348062 16718 348146 16954
rect 348382 16718 348414 16954
rect 347794 16634 348414 16718
rect 347794 16398 347826 16634
rect 348062 16398 348146 16634
rect 348382 16398 348414 16634
rect 383794 16718 383826 16954
rect 384062 16718 384146 16954
rect 384382 16718 384414 16954
rect 383794 16634 384414 16718
rect 383794 16398 383826 16634
rect 384062 16398 384146 16634
rect 384382 16398 384414 16634
rect 419794 16718 419826 16954
rect 420062 16718 420146 16954
rect 420382 16718 420414 16954
rect 419794 16634 420414 16718
rect 419794 16398 419826 16634
rect 420062 16398 420146 16634
rect 420382 16398 420414 16634
rect 455794 16718 455826 16954
rect 456062 16718 456146 16954
rect 456382 16718 456414 16954
rect 455794 16634 456414 16718
rect 455794 16398 455826 16634
rect 456062 16398 456146 16634
rect 456382 16398 456414 16634
rect 491794 16718 491826 16954
rect 492062 16718 492146 16954
rect 492382 16718 492414 16954
rect 491794 16634 492414 16718
rect 491794 16398 491826 16634
rect 492062 16398 492146 16634
rect 492382 16398 492414 16634
rect 527794 16718 527826 16954
rect 528062 16718 528146 16954
rect 528382 16718 528414 16954
rect 527794 16634 528414 16718
rect 527794 16398 527826 16634
rect 528062 16398 528146 16634
rect 528382 16398 528414 16634
rect 563794 16718 563826 16954
rect 564062 16718 564146 16954
rect 564382 16718 564414 16954
rect 563794 16634 564414 16718
rect 563794 16398 563826 16634
rect 564062 16398 564146 16634
rect 564382 16398 564414 16634
rect 582294 16718 582326 16954
rect 582562 16718 582646 16954
rect 582882 16718 582914 16954
rect 582294 16634 582914 16718
rect 582294 16398 582326 16634
rect 582562 16398 582646 16634
rect 582882 16398 582914 16634
rect -2006 12218 -1974 12454
rect -1738 12218 -1654 12454
rect -1418 12218 -1386 12454
rect -2006 12134 -1386 12218
rect -2006 11898 -1974 12134
rect -1738 11898 -1654 12134
rect -1418 11898 -1386 12134
rect 5794 12218 5826 12454
rect 6062 12218 6146 12454
rect 6382 12218 6414 12454
rect 5794 12134 6414 12218
rect 5794 11898 5826 12134
rect 6062 11898 6146 12134
rect 6382 11898 6414 12134
rect 41794 12218 41826 12454
rect 42062 12218 42146 12454
rect 42382 12218 42414 12454
rect 41794 12134 42414 12218
rect 41794 11898 41826 12134
rect 42062 11898 42146 12134
rect 42382 11898 42414 12134
rect 77794 12218 77826 12454
rect 78062 12218 78146 12454
rect 78382 12218 78414 12454
rect 77794 12134 78414 12218
rect 77794 11898 77826 12134
rect 78062 11898 78146 12134
rect 78382 11898 78414 12134
rect 113794 12218 113826 12454
rect 114062 12218 114146 12454
rect 114382 12218 114414 12454
rect 113794 12134 114414 12218
rect 113794 11898 113826 12134
rect 114062 11898 114146 12134
rect 114382 11898 114414 12134
rect 149794 12218 149826 12454
rect 150062 12218 150146 12454
rect 150382 12218 150414 12454
rect 149794 12134 150414 12218
rect 149794 11898 149826 12134
rect 150062 11898 150146 12134
rect 150382 11898 150414 12134
rect 185794 12218 185826 12454
rect 186062 12218 186146 12454
rect 186382 12218 186414 12454
rect 185794 12134 186414 12218
rect 185794 11898 185826 12134
rect 186062 11898 186146 12134
rect 186382 11898 186414 12134
rect 221794 12218 221826 12454
rect 222062 12218 222146 12454
rect 222382 12218 222414 12454
rect 221794 12134 222414 12218
rect 221794 11898 221826 12134
rect 222062 11898 222146 12134
rect 222382 11898 222414 12134
rect 257794 12218 257826 12454
rect 258062 12218 258146 12454
rect 258382 12218 258414 12454
rect 257794 12134 258414 12218
rect 257794 11898 257826 12134
rect 258062 11898 258146 12134
rect 258382 11898 258414 12134
rect 293794 12218 293826 12454
rect 294062 12218 294146 12454
rect 294382 12218 294414 12454
rect 293794 12134 294414 12218
rect 293794 11898 293826 12134
rect 294062 11898 294146 12134
rect 294382 11898 294414 12134
rect 329794 12218 329826 12454
rect 330062 12218 330146 12454
rect 330382 12218 330414 12454
rect 329794 12134 330414 12218
rect 329794 11898 329826 12134
rect 330062 11898 330146 12134
rect 330382 11898 330414 12134
rect 365794 12218 365826 12454
rect 366062 12218 366146 12454
rect 366382 12218 366414 12454
rect 365794 12134 366414 12218
rect 365794 11898 365826 12134
rect 366062 11898 366146 12134
rect 366382 11898 366414 12134
rect 401794 12218 401826 12454
rect 402062 12218 402146 12454
rect 402382 12218 402414 12454
rect 401794 12134 402414 12218
rect 401794 11898 401826 12134
rect 402062 11898 402146 12134
rect 402382 11898 402414 12134
rect 437794 12218 437826 12454
rect 438062 12218 438146 12454
rect 438382 12218 438414 12454
rect 437794 12134 438414 12218
rect 437794 11898 437826 12134
rect 438062 11898 438146 12134
rect 438382 11898 438414 12134
rect 473794 12218 473826 12454
rect 474062 12218 474146 12454
rect 474382 12218 474414 12454
rect 473794 12134 474414 12218
rect 473794 11898 473826 12134
rect 474062 11898 474146 12134
rect 474382 11898 474414 12134
rect 509794 12218 509826 12454
rect 510062 12218 510146 12454
rect 510382 12218 510414 12454
rect 509794 12134 510414 12218
rect 509794 11898 509826 12134
rect 510062 11898 510146 12134
rect 510382 11898 510414 12134
rect 545794 12218 545826 12454
rect 546062 12218 546146 12454
rect 546382 12218 546414 12454
rect 545794 12134 546414 12218
rect 545794 11898 545826 12134
rect 546062 11898 546146 12134
rect 546382 11898 546414 12134
rect -2006 -346 -1386 11898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect 582294 -1306 582914 16398
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 696454 585930 704282
rect 585310 696218 585342 696454
rect 585578 696218 585662 696454
rect 585898 696218 585930 696454
rect 585310 696134 585930 696218
rect 585310 695898 585342 696134
rect 585578 695898 585662 696134
rect 585898 695898 585930 696134
rect 585310 660454 585930 695898
rect 585310 660218 585342 660454
rect 585578 660218 585662 660454
rect 585898 660218 585930 660454
rect 585310 660134 585930 660218
rect 585310 659898 585342 660134
rect 585578 659898 585662 660134
rect 585898 659898 585930 660134
rect 585310 624454 585930 659898
rect 585310 624218 585342 624454
rect 585578 624218 585662 624454
rect 585898 624218 585930 624454
rect 585310 624134 585930 624218
rect 585310 623898 585342 624134
rect 585578 623898 585662 624134
rect 585898 623898 585930 624134
rect 585310 588454 585930 623898
rect 585310 588218 585342 588454
rect 585578 588218 585662 588454
rect 585898 588218 585930 588454
rect 585310 588134 585930 588218
rect 585310 587898 585342 588134
rect 585578 587898 585662 588134
rect 585898 587898 585930 588134
rect 585310 552454 585930 587898
rect 585310 552218 585342 552454
rect 585578 552218 585662 552454
rect 585898 552218 585930 552454
rect 585310 552134 585930 552218
rect 585310 551898 585342 552134
rect 585578 551898 585662 552134
rect 585898 551898 585930 552134
rect 585310 516454 585930 551898
rect 585310 516218 585342 516454
rect 585578 516218 585662 516454
rect 585898 516218 585930 516454
rect 585310 516134 585930 516218
rect 585310 515898 585342 516134
rect 585578 515898 585662 516134
rect 585898 515898 585930 516134
rect 585310 480454 585930 515898
rect 585310 480218 585342 480454
rect 585578 480218 585662 480454
rect 585898 480218 585930 480454
rect 585310 480134 585930 480218
rect 585310 479898 585342 480134
rect 585578 479898 585662 480134
rect 585898 479898 585930 480134
rect 585310 444454 585930 479898
rect 585310 444218 585342 444454
rect 585578 444218 585662 444454
rect 585898 444218 585930 444454
rect 585310 444134 585930 444218
rect 585310 443898 585342 444134
rect 585578 443898 585662 444134
rect 585898 443898 585930 444134
rect 585310 408454 585930 443898
rect 585310 408218 585342 408454
rect 585578 408218 585662 408454
rect 585898 408218 585930 408454
rect 585310 408134 585930 408218
rect 585310 407898 585342 408134
rect 585578 407898 585662 408134
rect 585898 407898 585930 408134
rect 585310 372454 585930 407898
rect 585310 372218 585342 372454
rect 585578 372218 585662 372454
rect 585898 372218 585930 372454
rect 585310 372134 585930 372218
rect 585310 371898 585342 372134
rect 585578 371898 585662 372134
rect 585898 371898 585930 372134
rect 585310 336454 585930 371898
rect 585310 336218 585342 336454
rect 585578 336218 585662 336454
rect 585898 336218 585930 336454
rect 585310 336134 585930 336218
rect 585310 335898 585342 336134
rect 585578 335898 585662 336134
rect 585898 335898 585930 336134
rect 585310 300454 585930 335898
rect 585310 300218 585342 300454
rect 585578 300218 585662 300454
rect 585898 300218 585930 300454
rect 585310 300134 585930 300218
rect 585310 299898 585342 300134
rect 585578 299898 585662 300134
rect 585898 299898 585930 300134
rect 585310 264454 585930 299898
rect 585310 264218 585342 264454
rect 585578 264218 585662 264454
rect 585898 264218 585930 264454
rect 585310 264134 585930 264218
rect 585310 263898 585342 264134
rect 585578 263898 585662 264134
rect 585898 263898 585930 264134
rect 585310 228454 585930 263898
rect 585310 228218 585342 228454
rect 585578 228218 585662 228454
rect 585898 228218 585930 228454
rect 585310 228134 585930 228218
rect 585310 227898 585342 228134
rect 585578 227898 585662 228134
rect 585898 227898 585930 228134
rect 585310 192454 585930 227898
rect 585310 192218 585342 192454
rect 585578 192218 585662 192454
rect 585898 192218 585930 192454
rect 585310 192134 585930 192218
rect 585310 191898 585342 192134
rect 585578 191898 585662 192134
rect 585898 191898 585930 192134
rect 585310 156454 585930 191898
rect 585310 156218 585342 156454
rect 585578 156218 585662 156454
rect 585898 156218 585930 156454
rect 585310 156134 585930 156218
rect 585310 155898 585342 156134
rect 585578 155898 585662 156134
rect 585898 155898 585930 156134
rect 585310 120454 585930 155898
rect 585310 120218 585342 120454
rect 585578 120218 585662 120454
rect 585898 120218 585930 120454
rect 585310 120134 585930 120218
rect 585310 119898 585342 120134
rect 585578 119898 585662 120134
rect 585898 119898 585930 120134
rect 585310 84454 585930 119898
rect 585310 84218 585342 84454
rect 585578 84218 585662 84454
rect 585898 84218 585930 84454
rect 585310 84134 585930 84218
rect 585310 83898 585342 84134
rect 585578 83898 585662 84134
rect 585898 83898 585930 84134
rect 585310 48454 585930 83898
rect 585310 48218 585342 48454
rect 585578 48218 585662 48454
rect 585898 48218 585930 48454
rect 585310 48134 585930 48218
rect 585310 47898 585342 48134
rect 585578 47898 585662 48134
rect 585898 47898 585930 48134
rect 585310 12454 585930 47898
rect 585310 12218 585342 12454
rect 585578 12218 585662 12454
rect 585898 12218 585930 12454
rect 585310 12134 585930 12218
rect 585310 11898 585342 12134
rect 585578 11898 585662 12134
rect 585898 11898 585930 12134
rect 585310 -346 585930 11898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 700954 586890 705242
rect 586270 700718 586302 700954
rect 586538 700718 586622 700954
rect 586858 700718 586890 700954
rect 586270 700634 586890 700718
rect 586270 700398 586302 700634
rect 586538 700398 586622 700634
rect 586858 700398 586890 700634
rect 586270 664954 586890 700398
rect 586270 664718 586302 664954
rect 586538 664718 586622 664954
rect 586858 664718 586890 664954
rect 586270 664634 586890 664718
rect 586270 664398 586302 664634
rect 586538 664398 586622 664634
rect 586858 664398 586890 664634
rect 586270 628954 586890 664398
rect 586270 628718 586302 628954
rect 586538 628718 586622 628954
rect 586858 628718 586890 628954
rect 586270 628634 586890 628718
rect 586270 628398 586302 628634
rect 586538 628398 586622 628634
rect 586858 628398 586890 628634
rect 586270 592954 586890 628398
rect 586270 592718 586302 592954
rect 586538 592718 586622 592954
rect 586858 592718 586890 592954
rect 586270 592634 586890 592718
rect 586270 592398 586302 592634
rect 586538 592398 586622 592634
rect 586858 592398 586890 592634
rect 586270 556954 586890 592398
rect 586270 556718 586302 556954
rect 586538 556718 586622 556954
rect 586858 556718 586890 556954
rect 586270 556634 586890 556718
rect 586270 556398 586302 556634
rect 586538 556398 586622 556634
rect 586858 556398 586890 556634
rect 586270 520954 586890 556398
rect 586270 520718 586302 520954
rect 586538 520718 586622 520954
rect 586858 520718 586890 520954
rect 586270 520634 586890 520718
rect 586270 520398 586302 520634
rect 586538 520398 586622 520634
rect 586858 520398 586890 520634
rect 586270 484954 586890 520398
rect 586270 484718 586302 484954
rect 586538 484718 586622 484954
rect 586858 484718 586890 484954
rect 586270 484634 586890 484718
rect 586270 484398 586302 484634
rect 586538 484398 586622 484634
rect 586858 484398 586890 484634
rect 586270 448954 586890 484398
rect 586270 448718 586302 448954
rect 586538 448718 586622 448954
rect 586858 448718 586890 448954
rect 586270 448634 586890 448718
rect 586270 448398 586302 448634
rect 586538 448398 586622 448634
rect 586858 448398 586890 448634
rect 586270 412954 586890 448398
rect 586270 412718 586302 412954
rect 586538 412718 586622 412954
rect 586858 412718 586890 412954
rect 586270 412634 586890 412718
rect 586270 412398 586302 412634
rect 586538 412398 586622 412634
rect 586858 412398 586890 412634
rect 586270 376954 586890 412398
rect 586270 376718 586302 376954
rect 586538 376718 586622 376954
rect 586858 376718 586890 376954
rect 586270 376634 586890 376718
rect 586270 376398 586302 376634
rect 586538 376398 586622 376634
rect 586858 376398 586890 376634
rect 586270 340954 586890 376398
rect 586270 340718 586302 340954
rect 586538 340718 586622 340954
rect 586858 340718 586890 340954
rect 586270 340634 586890 340718
rect 586270 340398 586302 340634
rect 586538 340398 586622 340634
rect 586858 340398 586890 340634
rect 586270 304954 586890 340398
rect 586270 304718 586302 304954
rect 586538 304718 586622 304954
rect 586858 304718 586890 304954
rect 586270 304634 586890 304718
rect 586270 304398 586302 304634
rect 586538 304398 586622 304634
rect 586858 304398 586890 304634
rect 586270 268954 586890 304398
rect 586270 268718 586302 268954
rect 586538 268718 586622 268954
rect 586858 268718 586890 268954
rect 586270 268634 586890 268718
rect 586270 268398 586302 268634
rect 586538 268398 586622 268634
rect 586858 268398 586890 268634
rect 586270 232954 586890 268398
rect 586270 232718 586302 232954
rect 586538 232718 586622 232954
rect 586858 232718 586890 232954
rect 586270 232634 586890 232718
rect 586270 232398 586302 232634
rect 586538 232398 586622 232634
rect 586858 232398 586890 232634
rect 586270 196954 586890 232398
rect 586270 196718 586302 196954
rect 586538 196718 586622 196954
rect 586858 196718 586890 196954
rect 586270 196634 586890 196718
rect 586270 196398 586302 196634
rect 586538 196398 586622 196634
rect 586858 196398 586890 196634
rect 586270 160954 586890 196398
rect 586270 160718 586302 160954
rect 586538 160718 586622 160954
rect 586858 160718 586890 160954
rect 586270 160634 586890 160718
rect 586270 160398 586302 160634
rect 586538 160398 586622 160634
rect 586858 160398 586890 160634
rect 586270 124954 586890 160398
rect 586270 124718 586302 124954
rect 586538 124718 586622 124954
rect 586858 124718 586890 124954
rect 586270 124634 586890 124718
rect 586270 124398 586302 124634
rect 586538 124398 586622 124634
rect 586858 124398 586890 124634
rect 586270 88954 586890 124398
rect 586270 88718 586302 88954
rect 586538 88718 586622 88954
rect 586858 88718 586890 88954
rect 586270 88634 586890 88718
rect 586270 88398 586302 88634
rect 586538 88398 586622 88634
rect 586858 88398 586890 88634
rect 586270 52954 586890 88398
rect 586270 52718 586302 52954
rect 586538 52718 586622 52954
rect 586858 52718 586890 52954
rect 586270 52634 586890 52718
rect 586270 52398 586302 52634
rect 586538 52398 586622 52634
rect 586858 52398 586890 52634
rect 586270 16954 586890 52398
rect 586270 16718 586302 16954
rect 586538 16718 586622 16954
rect 586858 16718 586890 16954
rect 586270 16634 586890 16718
rect 586270 16398 586302 16634
rect 586538 16398 586622 16634
rect 586858 16398 586890 16634
rect 582294 -1542 582326 -1306
rect 582562 -1542 582646 -1306
rect 582882 -1542 582914 -1306
rect 582294 -1626 582914 -1542
rect 582294 -1862 582326 -1626
rect 582562 -1862 582646 -1626
rect 582882 -1862 582914 -1626
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 582294 -7654 582914 -1862
rect 586270 -1306 586890 16398
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 -2266 587850 706202
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 -3226 588810 707162
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 -4186 589770 708122
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 -5146 590730 709082
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 -6106 591690 710042
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 -7066 592650 711002
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 582326 705562 582562 705798
rect 582646 705562 582882 705798
rect 582326 705242 582562 705478
rect 582646 705242 582882 705478
rect -2934 700718 -2698 700954
rect -2614 700718 -2378 700954
rect -2934 700398 -2698 700634
rect -2614 700398 -2378 700634
rect -2934 664718 -2698 664954
rect -2614 664718 -2378 664954
rect -2934 664398 -2698 664634
rect -2614 664398 -2378 664634
rect -2934 628718 -2698 628954
rect -2614 628718 -2378 628954
rect -2934 628398 -2698 628634
rect -2614 628398 -2378 628634
rect -2934 592718 -2698 592954
rect -2614 592718 -2378 592954
rect -2934 592398 -2698 592634
rect -2614 592398 -2378 592634
rect -2934 556718 -2698 556954
rect -2614 556718 -2378 556954
rect -2934 556398 -2698 556634
rect -2614 556398 -2378 556634
rect -2934 520718 -2698 520954
rect -2614 520718 -2378 520954
rect -2934 520398 -2698 520634
rect -2614 520398 -2378 520634
rect -2934 484718 -2698 484954
rect -2614 484718 -2378 484954
rect -2934 484398 -2698 484634
rect -2614 484398 -2378 484634
rect -2934 448718 -2698 448954
rect -2614 448718 -2378 448954
rect -2934 448398 -2698 448634
rect -2614 448398 -2378 448634
rect -2934 412718 -2698 412954
rect -2614 412718 -2378 412954
rect -2934 412398 -2698 412634
rect -2614 412398 -2378 412634
rect -2934 376718 -2698 376954
rect -2614 376718 -2378 376954
rect -2934 376398 -2698 376634
rect -2614 376398 -2378 376634
rect -2934 340718 -2698 340954
rect -2614 340718 -2378 340954
rect -2934 340398 -2698 340634
rect -2614 340398 -2378 340634
rect -2934 304718 -2698 304954
rect -2614 304718 -2378 304954
rect -2934 304398 -2698 304634
rect -2614 304398 -2378 304634
rect -2934 268718 -2698 268954
rect -2614 268718 -2378 268954
rect -2934 268398 -2698 268634
rect -2614 268398 -2378 268634
rect -2934 232718 -2698 232954
rect -2614 232718 -2378 232954
rect -2934 232398 -2698 232634
rect -2614 232398 -2378 232634
rect -2934 196718 -2698 196954
rect -2614 196718 -2378 196954
rect -2934 196398 -2698 196634
rect -2614 196398 -2378 196634
rect -2934 160718 -2698 160954
rect -2614 160718 -2378 160954
rect -2934 160398 -2698 160634
rect -2614 160398 -2378 160634
rect -2934 124718 -2698 124954
rect -2614 124718 -2378 124954
rect -2934 124398 -2698 124634
rect -2614 124398 -2378 124634
rect -2934 88718 -2698 88954
rect -2614 88718 -2378 88954
rect -2934 88398 -2698 88634
rect -2614 88398 -2378 88634
rect -2934 52718 -2698 52954
rect -2614 52718 -2378 52954
rect -2934 52398 -2698 52634
rect -2614 52398 -2378 52634
rect -2934 16718 -2698 16954
rect -2614 16718 -2378 16954
rect -2934 16398 -2698 16634
rect -2614 16398 -2378 16634
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 582326 700718 582562 700954
rect 582646 700718 582882 700954
rect 582326 700398 582562 700634
rect 582646 700398 582882 700634
rect -1974 696218 -1738 696454
rect -1654 696218 -1418 696454
rect -1974 695898 -1738 696134
rect -1654 695898 -1418 696134
rect 5826 696218 6062 696454
rect 6146 696218 6382 696454
rect 5826 695898 6062 696134
rect 6146 695898 6382 696134
rect 41826 696218 42062 696454
rect 42146 696218 42382 696454
rect 41826 695898 42062 696134
rect 42146 695898 42382 696134
rect 77826 696218 78062 696454
rect 78146 696218 78382 696454
rect 77826 695898 78062 696134
rect 78146 695898 78382 696134
rect 113826 696218 114062 696454
rect 114146 696218 114382 696454
rect 113826 695898 114062 696134
rect 114146 695898 114382 696134
rect 149826 696218 150062 696454
rect 150146 696218 150382 696454
rect 149826 695898 150062 696134
rect 150146 695898 150382 696134
rect 185826 696218 186062 696454
rect 186146 696218 186382 696454
rect 185826 695898 186062 696134
rect 186146 695898 186382 696134
rect 221826 696218 222062 696454
rect 222146 696218 222382 696454
rect 221826 695898 222062 696134
rect 222146 695898 222382 696134
rect 257826 696218 258062 696454
rect 258146 696218 258382 696454
rect 257826 695898 258062 696134
rect 258146 695898 258382 696134
rect 293826 696218 294062 696454
rect 294146 696218 294382 696454
rect 293826 695898 294062 696134
rect 294146 695898 294382 696134
rect 329826 696218 330062 696454
rect 330146 696218 330382 696454
rect 329826 695898 330062 696134
rect 330146 695898 330382 696134
rect 365826 696218 366062 696454
rect 366146 696218 366382 696454
rect 365826 695898 366062 696134
rect 366146 695898 366382 696134
rect 401826 696218 402062 696454
rect 402146 696218 402382 696454
rect 401826 695898 402062 696134
rect 402146 695898 402382 696134
rect 437826 696218 438062 696454
rect 438146 696218 438382 696454
rect 437826 695898 438062 696134
rect 438146 695898 438382 696134
rect 473826 696218 474062 696454
rect 474146 696218 474382 696454
rect 473826 695898 474062 696134
rect 474146 695898 474382 696134
rect 509826 696218 510062 696454
rect 510146 696218 510382 696454
rect 509826 695898 510062 696134
rect 510146 695898 510382 696134
rect 545826 696218 546062 696454
rect 546146 696218 546382 696454
rect 545826 695898 546062 696134
rect 546146 695898 546382 696134
rect 13198 664718 13434 664954
rect 13518 664718 13754 664954
rect 13198 664398 13434 664634
rect 13518 664398 13754 664634
rect 167826 664718 168062 664954
rect 168146 664718 168382 664954
rect 167826 664398 168062 664634
rect 168146 664398 168382 664634
rect 291590 664718 291826 664954
rect 291910 664718 292146 664954
rect 291590 664398 291826 664634
rect 291910 664398 292146 664634
rect 419826 664718 420062 664954
rect 420146 664718 420382 664954
rect 419826 664398 420062 664634
rect 420146 664398 420382 664634
rect 563826 664718 564062 664954
rect 564146 664718 564382 664954
rect 563826 664398 564062 664634
rect 564146 664398 564382 664634
rect 582326 664718 582562 664954
rect 582646 664718 582882 664954
rect 582326 664398 582562 664634
rect 582646 664398 582882 664634
rect -1974 660218 -1738 660454
rect -1654 660218 -1418 660454
rect -1974 659898 -1738 660134
rect -1654 659898 -1418 660134
rect 5826 660218 6062 660454
rect 6146 660218 6382 660454
rect 5826 659898 6062 660134
rect 6146 659898 6382 660134
rect 173094 660218 173330 660454
rect 173414 660218 173650 660454
rect 173094 659898 173330 660134
rect 173414 659898 173650 660134
rect 293826 660218 294062 660454
rect 294146 660218 294382 660454
rect 293826 659898 294062 660134
rect 294146 659898 294382 660134
rect 401826 660218 402062 660454
rect 402146 660218 402382 660454
rect 401826 659898 402062 660134
rect 402146 659898 402382 660134
rect 570350 660218 570586 660454
rect 570670 660218 570906 660454
rect 570350 659898 570586 660134
rect 570670 659898 570906 660134
rect 13198 628718 13434 628954
rect 13518 628718 13754 628954
rect 13198 628398 13434 628634
rect 13518 628398 13754 628634
rect 167826 628718 168062 628954
rect 168146 628718 168382 628954
rect 167826 628398 168062 628634
rect 168146 628398 168382 628634
rect 291590 628718 291826 628954
rect 291910 628718 292146 628954
rect 291590 628398 291826 628634
rect 291910 628398 292146 628634
rect 419826 628718 420062 628954
rect 420146 628718 420382 628954
rect 419826 628398 420062 628634
rect 420146 628398 420382 628634
rect 563826 628718 564062 628954
rect 564146 628718 564382 628954
rect 563826 628398 564062 628634
rect 564146 628398 564382 628634
rect 582326 628718 582562 628954
rect 582646 628718 582882 628954
rect 582326 628398 582562 628634
rect 582646 628398 582882 628634
rect -1974 624218 -1738 624454
rect -1654 624218 -1418 624454
rect -1974 623898 -1738 624134
rect -1654 623898 -1418 624134
rect 5826 624218 6062 624454
rect 6146 624218 6382 624454
rect 5826 623898 6062 624134
rect 6146 623898 6382 624134
rect 173094 624218 173330 624454
rect 173414 624218 173650 624454
rect 173094 623898 173330 624134
rect 173414 623898 173650 624134
rect 293826 624218 294062 624454
rect 294146 624218 294382 624454
rect 293826 623898 294062 624134
rect 294146 623898 294382 624134
rect 401826 624218 402062 624454
rect 402146 624218 402382 624454
rect 401826 623898 402062 624134
rect 402146 623898 402382 624134
rect 570350 624218 570586 624454
rect 570670 624218 570906 624454
rect 570350 623898 570586 624134
rect 570670 623898 570906 624134
rect 23826 592718 24062 592954
rect 24146 592718 24382 592954
rect 23826 592398 24062 592634
rect 24146 592398 24382 592634
rect 59826 592718 60062 592954
rect 60146 592718 60382 592954
rect 59826 592398 60062 592634
rect 60146 592398 60382 592634
rect 95826 592718 96062 592954
rect 96146 592718 96382 592954
rect 95826 592398 96062 592634
rect 96146 592398 96382 592634
rect 131826 592718 132062 592954
rect 132146 592718 132382 592954
rect 131826 592398 132062 592634
rect 132146 592398 132382 592634
rect 167826 592718 168062 592954
rect 168146 592718 168382 592954
rect 167826 592398 168062 592634
rect 168146 592398 168382 592634
rect 291590 592718 291826 592954
rect 291910 592718 292146 592954
rect 291590 592398 291826 592634
rect 291910 592398 292146 592634
rect 419826 592718 420062 592954
rect 420146 592718 420382 592954
rect 419826 592398 420062 592634
rect 420146 592398 420382 592634
rect 455826 592718 456062 592954
rect 456146 592718 456382 592954
rect 455826 592398 456062 592634
rect 456146 592398 456382 592634
rect 491826 592718 492062 592954
rect 492146 592718 492382 592954
rect 491826 592398 492062 592634
rect 492146 592398 492382 592634
rect 527826 592718 528062 592954
rect 528146 592718 528382 592954
rect 527826 592398 528062 592634
rect 528146 592398 528382 592634
rect 563826 592718 564062 592954
rect 564146 592718 564382 592954
rect 563826 592398 564062 592634
rect 564146 592398 564382 592634
rect 582326 592718 582562 592954
rect 582646 592718 582882 592954
rect 582326 592398 582562 592634
rect 582646 592398 582882 592634
rect -1974 588218 -1738 588454
rect -1654 588218 -1418 588454
rect -1974 587898 -1738 588134
rect -1654 587898 -1418 588134
rect 5826 588218 6062 588454
rect 6146 588218 6382 588454
rect 5826 587898 6062 588134
rect 6146 587898 6382 588134
rect 41826 588218 42062 588454
rect 42146 588218 42382 588454
rect 41826 587898 42062 588134
rect 42146 587898 42382 588134
rect 77826 588218 78062 588454
rect 78146 588218 78382 588454
rect 77826 587898 78062 588134
rect 78146 587898 78382 588134
rect 113826 588218 114062 588454
rect 114146 588218 114382 588454
rect 113826 587898 114062 588134
rect 114146 587898 114382 588134
rect 149826 588218 150062 588454
rect 150146 588218 150382 588454
rect 149826 587898 150062 588134
rect 150146 587898 150382 588134
rect 185826 588218 186062 588454
rect 186146 588218 186382 588454
rect 185826 587898 186062 588134
rect 186146 587898 186382 588134
rect 221826 588218 222062 588454
rect 222146 588218 222382 588454
rect 221826 587898 222062 588134
rect 222146 587898 222382 588134
rect 257826 588218 258062 588454
rect 258146 588218 258382 588454
rect 257826 587898 258062 588134
rect 258146 587898 258382 588134
rect 293826 588218 294062 588454
rect 294146 588218 294382 588454
rect 293826 587898 294062 588134
rect 294146 587898 294382 588134
rect 329826 588218 330062 588454
rect 330146 588218 330382 588454
rect 329826 587898 330062 588134
rect 330146 587898 330382 588134
rect 365826 588218 366062 588454
rect 366146 588218 366382 588454
rect 365826 587898 366062 588134
rect 366146 587898 366382 588134
rect 401826 588218 402062 588454
rect 402146 588218 402382 588454
rect 401826 587898 402062 588134
rect 402146 587898 402382 588134
rect 437826 588218 438062 588454
rect 438146 588218 438382 588454
rect 437826 587898 438062 588134
rect 438146 587898 438382 588134
rect 473826 588218 474062 588454
rect 474146 588218 474382 588454
rect 473826 587898 474062 588134
rect 474146 587898 474382 588134
rect 509826 588218 510062 588454
rect 510146 588218 510382 588454
rect 509826 587898 510062 588134
rect 510146 587898 510382 588134
rect 545826 588218 546062 588454
rect 546146 588218 546382 588454
rect 545826 587898 546062 588134
rect 546146 587898 546382 588134
rect 13198 556718 13434 556954
rect 13518 556718 13754 556954
rect 13198 556398 13434 556634
rect 13518 556398 13754 556634
rect 167826 556718 168062 556954
rect 168146 556718 168382 556954
rect 167826 556398 168062 556634
rect 168146 556398 168382 556634
rect 203826 556718 204062 556954
rect 204146 556718 204382 556954
rect 203826 556398 204062 556634
rect 204146 556398 204382 556634
rect 239826 556718 240062 556954
rect 240146 556718 240382 556954
rect 239826 556398 240062 556634
rect 240146 556398 240382 556634
rect 275826 556718 276062 556954
rect 276146 556718 276382 556954
rect 275826 556398 276062 556634
rect 276146 556398 276382 556634
rect 311826 556718 312062 556954
rect 312146 556718 312382 556954
rect 311826 556398 312062 556634
rect 312146 556398 312382 556634
rect 347826 556718 348062 556954
rect 348146 556718 348382 556954
rect 347826 556398 348062 556634
rect 348146 556398 348382 556634
rect 383826 556718 384062 556954
rect 384146 556718 384382 556954
rect 383826 556398 384062 556634
rect 384146 556398 384382 556634
rect 419826 556718 420062 556954
rect 420146 556718 420382 556954
rect 419826 556398 420062 556634
rect 420146 556398 420382 556634
rect 563826 556718 564062 556954
rect 564146 556718 564382 556954
rect 563826 556398 564062 556634
rect 564146 556398 564382 556634
rect 582326 556718 582562 556954
rect 582646 556718 582882 556954
rect 582326 556398 582562 556634
rect 582646 556398 582882 556634
rect -1974 552218 -1738 552454
rect -1654 552218 -1418 552454
rect -1974 551898 -1738 552134
rect -1654 551898 -1418 552134
rect 5826 552218 6062 552454
rect 6146 552218 6382 552454
rect 5826 551898 6062 552134
rect 6146 551898 6382 552134
rect 185826 552218 186062 552454
rect 186146 552218 186382 552454
rect 185826 551898 186062 552134
rect 186146 551898 186382 552134
rect 221826 552218 222062 552454
rect 222146 552218 222382 552454
rect 221826 551898 222062 552134
rect 222146 551898 222382 552134
rect 257826 552218 258062 552454
rect 258146 552218 258382 552454
rect 257826 551898 258062 552134
rect 258146 551898 258382 552134
rect 293826 552218 294062 552454
rect 294146 552218 294382 552454
rect 293826 551898 294062 552134
rect 294146 551898 294382 552134
rect 329826 552218 330062 552454
rect 330146 552218 330382 552454
rect 329826 551898 330062 552134
rect 330146 551898 330382 552134
rect 365826 552218 366062 552454
rect 366146 552218 366382 552454
rect 365826 551898 366062 552134
rect 366146 551898 366382 552134
rect 401826 552218 402062 552454
rect 402146 552218 402382 552454
rect 401826 551898 402062 552134
rect 402146 551898 402382 552134
rect 570350 552218 570586 552454
rect 570670 552218 570906 552454
rect 570350 551898 570586 552134
rect 570670 551898 570906 552134
rect 13198 520718 13434 520954
rect 13518 520718 13754 520954
rect 13198 520398 13434 520634
rect 13518 520398 13754 520634
rect 167826 520718 168062 520954
rect 168146 520718 168382 520954
rect 167826 520398 168062 520634
rect 168146 520398 168382 520634
rect 203826 520718 204062 520954
rect 204146 520718 204382 520954
rect 203826 520398 204062 520634
rect 204146 520398 204382 520634
rect 239826 520718 240062 520954
rect 240146 520718 240382 520954
rect 239826 520398 240062 520634
rect 240146 520398 240382 520634
rect 275826 520718 276062 520954
rect 276146 520718 276382 520954
rect 275826 520398 276062 520634
rect 276146 520398 276382 520634
rect 311826 520718 312062 520954
rect 312146 520718 312382 520954
rect 311826 520398 312062 520634
rect 312146 520398 312382 520634
rect 347826 520718 348062 520954
rect 348146 520718 348382 520954
rect 347826 520398 348062 520634
rect 348146 520398 348382 520634
rect 383826 520718 384062 520954
rect 384146 520718 384382 520954
rect 383826 520398 384062 520634
rect 384146 520398 384382 520634
rect 419826 520718 420062 520954
rect 420146 520718 420382 520954
rect 419826 520398 420062 520634
rect 420146 520398 420382 520634
rect 563826 520718 564062 520954
rect 564146 520718 564382 520954
rect 563826 520398 564062 520634
rect 564146 520398 564382 520634
rect 582326 520718 582562 520954
rect 582646 520718 582882 520954
rect 582326 520398 582562 520634
rect 582646 520398 582882 520634
rect -1974 516218 -1738 516454
rect -1654 516218 -1418 516454
rect -1974 515898 -1738 516134
rect -1654 515898 -1418 516134
rect 5826 516218 6062 516454
rect 6146 516218 6382 516454
rect 5826 515898 6062 516134
rect 6146 515898 6382 516134
rect 185826 516218 186062 516454
rect 186146 516218 186382 516454
rect 185826 515898 186062 516134
rect 186146 515898 186382 516134
rect 221826 516218 222062 516454
rect 222146 516218 222382 516454
rect 221826 515898 222062 516134
rect 222146 515898 222382 516134
rect 257826 516218 258062 516454
rect 258146 516218 258382 516454
rect 257826 515898 258062 516134
rect 258146 515898 258382 516134
rect 293826 516218 294062 516454
rect 294146 516218 294382 516454
rect 293826 515898 294062 516134
rect 294146 515898 294382 516134
rect 329826 516218 330062 516454
rect 330146 516218 330382 516454
rect 329826 515898 330062 516134
rect 330146 515898 330382 516134
rect 365826 516218 366062 516454
rect 366146 516218 366382 516454
rect 365826 515898 366062 516134
rect 366146 515898 366382 516134
rect 401826 516218 402062 516454
rect 402146 516218 402382 516454
rect 401826 515898 402062 516134
rect 402146 515898 402382 516134
rect 570350 516218 570586 516454
rect 570670 516218 570906 516454
rect 570350 515898 570586 516134
rect 570670 515898 570906 516134
rect 23826 484718 24062 484954
rect 24146 484718 24382 484954
rect 23826 484398 24062 484634
rect 24146 484398 24382 484634
rect 59826 484718 60062 484954
rect 60146 484718 60382 484954
rect 59826 484398 60062 484634
rect 60146 484398 60382 484634
rect 95826 484718 96062 484954
rect 96146 484718 96382 484954
rect 95826 484398 96062 484634
rect 96146 484398 96382 484634
rect 131826 484718 132062 484954
rect 132146 484718 132382 484954
rect 131826 484398 132062 484634
rect 132146 484398 132382 484634
rect 167826 484718 168062 484954
rect 168146 484718 168382 484954
rect 167826 484398 168062 484634
rect 168146 484398 168382 484634
rect 203826 484718 204062 484954
rect 204146 484718 204382 484954
rect 203826 484398 204062 484634
rect 204146 484398 204382 484634
rect 239826 484718 240062 484954
rect 240146 484718 240382 484954
rect 239826 484398 240062 484634
rect 240146 484398 240382 484634
rect 275826 484718 276062 484954
rect 276146 484718 276382 484954
rect 275826 484398 276062 484634
rect 276146 484398 276382 484634
rect 311826 484718 312062 484954
rect 312146 484718 312382 484954
rect 311826 484398 312062 484634
rect 312146 484398 312382 484634
rect 347826 484718 348062 484954
rect 348146 484718 348382 484954
rect 347826 484398 348062 484634
rect 348146 484398 348382 484634
rect 383826 484718 384062 484954
rect 384146 484718 384382 484954
rect 383826 484398 384062 484634
rect 384146 484398 384382 484634
rect 419826 484718 420062 484954
rect 420146 484718 420382 484954
rect 419826 484398 420062 484634
rect 420146 484398 420382 484634
rect 455826 484718 456062 484954
rect 456146 484718 456382 484954
rect 455826 484398 456062 484634
rect 456146 484398 456382 484634
rect 491826 484718 492062 484954
rect 492146 484718 492382 484954
rect 491826 484398 492062 484634
rect 492146 484398 492382 484634
rect 527826 484718 528062 484954
rect 528146 484718 528382 484954
rect 527826 484398 528062 484634
rect 528146 484398 528382 484634
rect 563826 484718 564062 484954
rect 564146 484718 564382 484954
rect 563826 484398 564062 484634
rect 564146 484398 564382 484634
rect 582326 484718 582562 484954
rect 582646 484718 582882 484954
rect 582326 484398 582562 484634
rect 582646 484398 582882 484634
rect -1974 480218 -1738 480454
rect -1654 480218 -1418 480454
rect -1974 479898 -1738 480134
rect -1654 479898 -1418 480134
rect 5826 480218 6062 480454
rect 6146 480218 6382 480454
rect 5826 479898 6062 480134
rect 6146 479898 6382 480134
rect 41826 480218 42062 480454
rect 42146 480218 42382 480454
rect 41826 479898 42062 480134
rect 42146 479898 42382 480134
rect 77826 480218 78062 480454
rect 78146 480218 78382 480454
rect 77826 479898 78062 480134
rect 78146 479898 78382 480134
rect 113826 480218 114062 480454
rect 114146 480218 114382 480454
rect 113826 479898 114062 480134
rect 114146 479898 114382 480134
rect 149826 480218 150062 480454
rect 150146 480218 150382 480454
rect 149826 479898 150062 480134
rect 150146 479898 150382 480134
rect 185826 480218 186062 480454
rect 186146 480218 186382 480454
rect 185826 479898 186062 480134
rect 186146 479898 186382 480134
rect 221826 480218 222062 480454
rect 222146 480218 222382 480454
rect 221826 479898 222062 480134
rect 222146 479898 222382 480134
rect 257826 480218 258062 480454
rect 258146 480218 258382 480454
rect 257826 479898 258062 480134
rect 258146 479898 258382 480134
rect 293826 480218 294062 480454
rect 294146 480218 294382 480454
rect 293826 479898 294062 480134
rect 294146 479898 294382 480134
rect 329826 480218 330062 480454
rect 330146 480218 330382 480454
rect 329826 479898 330062 480134
rect 330146 479898 330382 480134
rect 365826 480218 366062 480454
rect 366146 480218 366382 480454
rect 365826 479898 366062 480134
rect 366146 479898 366382 480134
rect 401826 480218 402062 480454
rect 402146 480218 402382 480454
rect 401826 479898 402062 480134
rect 402146 479898 402382 480134
rect 437826 480218 438062 480454
rect 438146 480218 438382 480454
rect 437826 479898 438062 480134
rect 438146 479898 438382 480134
rect 473826 480218 474062 480454
rect 474146 480218 474382 480454
rect 473826 479898 474062 480134
rect 474146 479898 474382 480134
rect 509826 480218 510062 480454
rect 510146 480218 510382 480454
rect 509826 479898 510062 480134
rect 510146 479898 510382 480134
rect 545826 480218 546062 480454
rect 546146 480218 546382 480454
rect 545826 479898 546062 480134
rect 546146 479898 546382 480134
rect 13198 448718 13434 448954
rect 13518 448718 13754 448954
rect 13198 448398 13434 448634
rect 13518 448398 13754 448634
rect 167826 448718 168062 448954
rect 168146 448718 168382 448954
rect 167826 448398 168062 448634
rect 168146 448398 168382 448634
rect 203826 448718 204062 448954
rect 204146 448718 204382 448954
rect 203826 448398 204062 448634
rect 204146 448398 204382 448634
rect 239826 448718 240062 448954
rect 240146 448718 240382 448954
rect 239826 448398 240062 448634
rect 240146 448398 240382 448634
rect 275826 448718 276062 448954
rect 276146 448718 276382 448954
rect 275826 448398 276062 448634
rect 276146 448398 276382 448634
rect 311826 448718 312062 448954
rect 312146 448718 312382 448954
rect 311826 448398 312062 448634
rect 312146 448398 312382 448634
rect 347826 448718 348062 448954
rect 348146 448718 348382 448954
rect 347826 448398 348062 448634
rect 348146 448398 348382 448634
rect 383826 448718 384062 448954
rect 384146 448718 384382 448954
rect 383826 448398 384062 448634
rect 384146 448398 384382 448634
rect 419826 448718 420062 448954
rect 420146 448718 420382 448954
rect 419826 448398 420062 448634
rect 420146 448398 420382 448634
rect 563826 448718 564062 448954
rect 564146 448718 564382 448954
rect 563826 448398 564062 448634
rect 564146 448398 564382 448634
rect 582326 448718 582562 448954
rect 582646 448718 582882 448954
rect 582326 448398 582562 448634
rect 582646 448398 582882 448634
rect -1974 444218 -1738 444454
rect -1654 444218 -1418 444454
rect -1974 443898 -1738 444134
rect -1654 443898 -1418 444134
rect 5826 444218 6062 444454
rect 6146 444218 6382 444454
rect 5826 443898 6062 444134
rect 6146 443898 6382 444134
rect 185826 444218 186062 444454
rect 186146 444218 186382 444454
rect 185826 443898 186062 444134
rect 186146 443898 186382 444134
rect 221826 444218 222062 444454
rect 222146 444218 222382 444454
rect 221826 443898 222062 444134
rect 222146 443898 222382 444134
rect 257826 444218 258062 444454
rect 258146 444218 258382 444454
rect 257826 443898 258062 444134
rect 258146 443898 258382 444134
rect 293826 444218 294062 444454
rect 294146 444218 294382 444454
rect 293826 443898 294062 444134
rect 294146 443898 294382 444134
rect 329826 444218 330062 444454
rect 330146 444218 330382 444454
rect 329826 443898 330062 444134
rect 330146 443898 330382 444134
rect 365826 444218 366062 444454
rect 366146 444218 366382 444454
rect 365826 443898 366062 444134
rect 366146 443898 366382 444134
rect 401826 444218 402062 444454
rect 402146 444218 402382 444454
rect 401826 443898 402062 444134
rect 402146 443898 402382 444134
rect 570350 444218 570586 444454
rect 570670 444218 570906 444454
rect 570350 443898 570586 444134
rect 570670 443898 570906 444134
rect 13198 412718 13434 412954
rect 13518 412718 13754 412954
rect 13198 412398 13434 412634
rect 13518 412398 13754 412634
rect 167826 412718 168062 412954
rect 168146 412718 168382 412954
rect 167826 412398 168062 412634
rect 168146 412398 168382 412634
rect 203826 412718 204062 412954
rect 204146 412718 204382 412954
rect 203826 412398 204062 412634
rect 204146 412398 204382 412634
rect 239826 412718 240062 412954
rect 240146 412718 240382 412954
rect 239826 412398 240062 412634
rect 240146 412398 240382 412634
rect 275826 412718 276062 412954
rect 276146 412718 276382 412954
rect 275826 412398 276062 412634
rect 276146 412398 276382 412634
rect 311826 412718 312062 412954
rect 312146 412718 312382 412954
rect 311826 412398 312062 412634
rect 312146 412398 312382 412634
rect 347826 412718 348062 412954
rect 348146 412718 348382 412954
rect 347826 412398 348062 412634
rect 348146 412398 348382 412634
rect 383826 412718 384062 412954
rect 384146 412718 384382 412954
rect 383826 412398 384062 412634
rect 384146 412398 384382 412634
rect 419826 412718 420062 412954
rect 420146 412718 420382 412954
rect 419826 412398 420062 412634
rect 420146 412398 420382 412634
rect 563826 412718 564062 412954
rect 564146 412718 564382 412954
rect 563826 412398 564062 412634
rect 564146 412398 564382 412634
rect 582326 412718 582562 412954
rect 582646 412718 582882 412954
rect 582326 412398 582562 412634
rect 582646 412398 582882 412634
rect -1974 408218 -1738 408454
rect -1654 408218 -1418 408454
rect -1974 407898 -1738 408134
rect -1654 407898 -1418 408134
rect 5826 408218 6062 408454
rect 6146 408218 6382 408454
rect 5826 407898 6062 408134
rect 6146 407898 6382 408134
rect 185826 408218 186062 408454
rect 186146 408218 186382 408454
rect 185826 407898 186062 408134
rect 186146 407898 186382 408134
rect 221826 408218 222062 408454
rect 222146 408218 222382 408454
rect 221826 407898 222062 408134
rect 222146 407898 222382 408134
rect 257826 408218 258062 408454
rect 258146 408218 258382 408454
rect 257826 407898 258062 408134
rect 258146 407898 258382 408134
rect 293826 408218 294062 408454
rect 294146 408218 294382 408454
rect 293826 407898 294062 408134
rect 294146 407898 294382 408134
rect 329826 408218 330062 408454
rect 330146 408218 330382 408454
rect 329826 407898 330062 408134
rect 330146 407898 330382 408134
rect 365826 408218 366062 408454
rect 366146 408218 366382 408454
rect 365826 407898 366062 408134
rect 366146 407898 366382 408134
rect 401826 408218 402062 408454
rect 402146 408218 402382 408454
rect 401826 407898 402062 408134
rect 402146 407898 402382 408134
rect 570350 408218 570586 408454
rect 570670 408218 570906 408454
rect 570350 407898 570586 408134
rect 570670 407898 570906 408134
rect 13198 376718 13434 376954
rect 13518 376718 13754 376954
rect 13198 376398 13434 376634
rect 13518 376398 13754 376634
rect 167826 376718 168062 376954
rect 168146 376718 168382 376954
rect 167826 376398 168062 376634
rect 168146 376398 168382 376634
rect 203826 376718 204062 376954
rect 204146 376718 204382 376954
rect 203826 376398 204062 376634
rect 204146 376398 204382 376634
rect 239826 376718 240062 376954
rect 240146 376718 240382 376954
rect 239826 376398 240062 376634
rect 240146 376398 240382 376634
rect 275826 376718 276062 376954
rect 276146 376718 276382 376954
rect 275826 376398 276062 376634
rect 276146 376398 276382 376634
rect 311826 376718 312062 376954
rect 312146 376718 312382 376954
rect 311826 376398 312062 376634
rect 312146 376398 312382 376634
rect 347826 376718 348062 376954
rect 348146 376718 348382 376954
rect 347826 376398 348062 376634
rect 348146 376398 348382 376634
rect 383826 376718 384062 376954
rect 384146 376718 384382 376954
rect 383826 376398 384062 376634
rect 384146 376398 384382 376634
rect 419826 376718 420062 376954
rect 420146 376718 420382 376954
rect 419826 376398 420062 376634
rect 420146 376398 420382 376634
rect 563826 376718 564062 376954
rect 564146 376718 564382 376954
rect 563826 376398 564062 376634
rect 564146 376398 564382 376634
rect 582326 376718 582562 376954
rect 582646 376718 582882 376954
rect 582326 376398 582562 376634
rect 582646 376398 582882 376634
rect -1974 372218 -1738 372454
rect -1654 372218 -1418 372454
rect -1974 371898 -1738 372134
rect -1654 371898 -1418 372134
rect 5826 372218 6062 372454
rect 6146 372218 6382 372454
rect 5826 371898 6062 372134
rect 6146 371898 6382 372134
rect 185826 372218 186062 372454
rect 186146 372218 186382 372454
rect 185826 371898 186062 372134
rect 186146 371898 186382 372134
rect 221826 372218 222062 372454
rect 222146 372218 222382 372454
rect 221826 371898 222062 372134
rect 222146 371898 222382 372134
rect 257826 372218 258062 372454
rect 258146 372218 258382 372454
rect 257826 371898 258062 372134
rect 258146 371898 258382 372134
rect 293826 372218 294062 372454
rect 294146 372218 294382 372454
rect 293826 371898 294062 372134
rect 294146 371898 294382 372134
rect 329826 372218 330062 372454
rect 330146 372218 330382 372454
rect 329826 371898 330062 372134
rect 330146 371898 330382 372134
rect 365826 372218 366062 372454
rect 366146 372218 366382 372454
rect 365826 371898 366062 372134
rect 366146 371898 366382 372134
rect 401826 372218 402062 372454
rect 402146 372218 402382 372454
rect 401826 371898 402062 372134
rect 402146 371898 402382 372134
rect 570350 372218 570586 372454
rect 570670 372218 570906 372454
rect 570350 371898 570586 372134
rect 570670 371898 570906 372134
rect 13198 340718 13434 340954
rect 13518 340718 13754 340954
rect 13198 340398 13434 340634
rect 13518 340398 13754 340634
rect 167826 340718 168062 340954
rect 168146 340718 168382 340954
rect 167826 340398 168062 340634
rect 168146 340398 168382 340634
rect 203826 340718 204062 340954
rect 204146 340718 204382 340954
rect 203826 340398 204062 340634
rect 204146 340398 204382 340634
rect 239826 340718 240062 340954
rect 240146 340718 240382 340954
rect 239826 340398 240062 340634
rect 240146 340398 240382 340634
rect 275826 340718 276062 340954
rect 276146 340718 276382 340954
rect 275826 340398 276062 340634
rect 276146 340398 276382 340634
rect 311826 340718 312062 340954
rect 312146 340718 312382 340954
rect 311826 340398 312062 340634
rect 312146 340398 312382 340634
rect 347826 340718 348062 340954
rect 348146 340718 348382 340954
rect 347826 340398 348062 340634
rect 348146 340398 348382 340634
rect 383826 340718 384062 340954
rect 384146 340718 384382 340954
rect 383826 340398 384062 340634
rect 384146 340398 384382 340634
rect 419826 340718 420062 340954
rect 420146 340718 420382 340954
rect 419826 340398 420062 340634
rect 420146 340398 420382 340634
rect 563826 340718 564062 340954
rect 564146 340718 564382 340954
rect 563826 340398 564062 340634
rect 564146 340398 564382 340634
rect 582326 340718 582562 340954
rect 582646 340718 582882 340954
rect 582326 340398 582562 340634
rect 582646 340398 582882 340634
rect -1974 336218 -1738 336454
rect -1654 336218 -1418 336454
rect -1974 335898 -1738 336134
rect -1654 335898 -1418 336134
rect 5826 336218 6062 336454
rect 6146 336218 6382 336454
rect 5826 335898 6062 336134
rect 6146 335898 6382 336134
rect 185826 336218 186062 336454
rect 186146 336218 186382 336454
rect 185826 335898 186062 336134
rect 186146 335898 186382 336134
rect 221826 336218 222062 336454
rect 222146 336218 222382 336454
rect 221826 335898 222062 336134
rect 222146 335898 222382 336134
rect 257826 336218 258062 336454
rect 258146 336218 258382 336454
rect 257826 335898 258062 336134
rect 258146 335898 258382 336134
rect 293826 336218 294062 336454
rect 294146 336218 294382 336454
rect 293826 335898 294062 336134
rect 294146 335898 294382 336134
rect 329826 336218 330062 336454
rect 330146 336218 330382 336454
rect 329826 335898 330062 336134
rect 330146 335898 330382 336134
rect 365826 336218 366062 336454
rect 366146 336218 366382 336454
rect 365826 335898 366062 336134
rect 366146 335898 366382 336134
rect 401826 336218 402062 336454
rect 402146 336218 402382 336454
rect 401826 335898 402062 336134
rect 402146 335898 402382 336134
rect 570350 336218 570586 336454
rect 570670 336218 570906 336454
rect 570350 335898 570586 336134
rect 570670 335898 570906 336134
rect 13198 304718 13434 304954
rect 13518 304718 13754 304954
rect 13198 304398 13434 304634
rect 13518 304398 13754 304634
rect 167826 304718 168062 304954
rect 168146 304718 168382 304954
rect 167826 304398 168062 304634
rect 168146 304398 168382 304634
rect 203826 304718 204062 304954
rect 204146 304718 204382 304954
rect 203826 304398 204062 304634
rect 204146 304398 204382 304634
rect 239826 304718 240062 304954
rect 240146 304718 240382 304954
rect 239826 304398 240062 304634
rect 240146 304398 240382 304634
rect 275826 304718 276062 304954
rect 276146 304718 276382 304954
rect 275826 304398 276062 304634
rect 276146 304398 276382 304634
rect 311826 304718 312062 304954
rect 312146 304718 312382 304954
rect 311826 304398 312062 304634
rect 312146 304398 312382 304634
rect 347826 304718 348062 304954
rect 348146 304718 348382 304954
rect 347826 304398 348062 304634
rect 348146 304398 348382 304634
rect 383826 304718 384062 304954
rect 384146 304718 384382 304954
rect 383826 304398 384062 304634
rect 384146 304398 384382 304634
rect 419826 304718 420062 304954
rect 420146 304718 420382 304954
rect 419826 304398 420062 304634
rect 420146 304398 420382 304634
rect 563826 304718 564062 304954
rect 564146 304718 564382 304954
rect 563826 304398 564062 304634
rect 564146 304398 564382 304634
rect 582326 304718 582562 304954
rect 582646 304718 582882 304954
rect 582326 304398 582562 304634
rect 582646 304398 582882 304634
rect -1974 300218 -1738 300454
rect -1654 300218 -1418 300454
rect -1974 299898 -1738 300134
rect -1654 299898 -1418 300134
rect 5826 300218 6062 300454
rect 6146 300218 6382 300454
rect 5826 299898 6062 300134
rect 6146 299898 6382 300134
rect 185826 300218 186062 300454
rect 186146 300218 186382 300454
rect 185826 299898 186062 300134
rect 186146 299898 186382 300134
rect 221826 300218 222062 300454
rect 222146 300218 222382 300454
rect 221826 299898 222062 300134
rect 222146 299898 222382 300134
rect 257826 300218 258062 300454
rect 258146 300218 258382 300454
rect 257826 299898 258062 300134
rect 258146 299898 258382 300134
rect 293826 300218 294062 300454
rect 294146 300218 294382 300454
rect 293826 299898 294062 300134
rect 294146 299898 294382 300134
rect 329826 300218 330062 300454
rect 330146 300218 330382 300454
rect 329826 299898 330062 300134
rect 330146 299898 330382 300134
rect 365826 300218 366062 300454
rect 366146 300218 366382 300454
rect 365826 299898 366062 300134
rect 366146 299898 366382 300134
rect 401826 300218 402062 300454
rect 402146 300218 402382 300454
rect 401826 299898 402062 300134
rect 402146 299898 402382 300134
rect 570350 300218 570586 300454
rect 570670 300218 570906 300454
rect 570350 299898 570586 300134
rect 570670 299898 570906 300134
rect 13198 268718 13434 268954
rect 13518 268718 13754 268954
rect 13198 268398 13434 268634
rect 13518 268398 13754 268634
rect 167826 268718 168062 268954
rect 168146 268718 168382 268954
rect 167826 268398 168062 268634
rect 168146 268398 168382 268634
rect 203826 268718 204062 268954
rect 204146 268718 204382 268954
rect 203826 268398 204062 268634
rect 204146 268398 204382 268634
rect 239826 268718 240062 268954
rect 240146 268718 240382 268954
rect 239826 268398 240062 268634
rect 240146 268398 240382 268634
rect 275826 268718 276062 268954
rect 276146 268718 276382 268954
rect 275826 268398 276062 268634
rect 276146 268398 276382 268634
rect 311826 268718 312062 268954
rect 312146 268718 312382 268954
rect 311826 268398 312062 268634
rect 312146 268398 312382 268634
rect 347826 268718 348062 268954
rect 348146 268718 348382 268954
rect 347826 268398 348062 268634
rect 348146 268398 348382 268634
rect 383826 268718 384062 268954
rect 384146 268718 384382 268954
rect 383826 268398 384062 268634
rect 384146 268398 384382 268634
rect 419826 268718 420062 268954
rect 420146 268718 420382 268954
rect 419826 268398 420062 268634
rect 420146 268398 420382 268634
rect 563826 268718 564062 268954
rect 564146 268718 564382 268954
rect 563826 268398 564062 268634
rect 564146 268398 564382 268634
rect 582326 268718 582562 268954
rect 582646 268718 582882 268954
rect 582326 268398 582562 268634
rect 582646 268398 582882 268634
rect -1974 264218 -1738 264454
rect -1654 264218 -1418 264454
rect -1974 263898 -1738 264134
rect -1654 263898 -1418 264134
rect 5826 264218 6062 264454
rect 6146 264218 6382 264454
rect 5826 263898 6062 264134
rect 6146 263898 6382 264134
rect 185826 264218 186062 264454
rect 186146 264218 186382 264454
rect 185826 263898 186062 264134
rect 186146 263898 186382 264134
rect 221826 264218 222062 264454
rect 222146 264218 222382 264454
rect 221826 263898 222062 264134
rect 222146 263898 222382 264134
rect 257826 264218 258062 264454
rect 258146 264218 258382 264454
rect 257826 263898 258062 264134
rect 258146 263898 258382 264134
rect 293826 264218 294062 264454
rect 294146 264218 294382 264454
rect 293826 263898 294062 264134
rect 294146 263898 294382 264134
rect 329826 264218 330062 264454
rect 330146 264218 330382 264454
rect 329826 263898 330062 264134
rect 330146 263898 330382 264134
rect 365826 264218 366062 264454
rect 366146 264218 366382 264454
rect 365826 263898 366062 264134
rect 366146 263898 366382 264134
rect 401826 264218 402062 264454
rect 402146 264218 402382 264454
rect 401826 263898 402062 264134
rect 402146 263898 402382 264134
rect 570350 264218 570586 264454
rect 570670 264218 570906 264454
rect 570350 263898 570586 264134
rect 570670 263898 570906 264134
rect 23826 232718 24062 232954
rect 24146 232718 24382 232954
rect 23826 232398 24062 232634
rect 24146 232398 24382 232634
rect 59826 232718 60062 232954
rect 60146 232718 60382 232954
rect 59826 232398 60062 232634
rect 60146 232398 60382 232634
rect 95826 232718 96062 232954
rect 96146 232718 96382 232954
rect 95826 232398 96062 232634
rect 96146 232398 96382 232634
rect 131826 232718 132062 232954
rect 132146 232718 132382 232954
rect 131826 232398 132062 232634
rect 132146 232398 132382 232634
rect 167826 232718 168062 232954
rect 168146 232718 168382 232954
rect 167826 232398 168062 232634
rect 168146 232398 168382 232634
rect 203826 232718 204062 232954
rect 204146 232718 204382 232954
rect 203826 232398 204062 232634
rect 204146 232398 204382 232634
rect 239826 232718 240062 232954
rect 240146 232718 240382 232954
rect 239826 232398 240062 232634
rect 240146 232398 240382 232634
rect 275826 232718 276062 232954
rect 276146 232718 276382 232954
rect 275826 232398 276062 232634
rect 276146 232398 276382 232634
rect 311826 232718 312062 232954
rect 312146 232718 312382 232954
rect 311826 232398 312062 232634
rect 312146 232398 312382 232634
rect 347826 232718 348062 232954
rect 348146 232718 348382 232954
rect 347826 232398 348062 232634
rect 348146 232398 348382 232634
rect 383826 232718 384062 232954
rect 384146 232718 384382 232954
rect 383826 232398 384062 232634
rect 384146 232398 384382 232634
rect 419826 232718 420062 232954
rect 420146 232718 420382 232954
rect 419826 232398 420062 232634
rect 420146 232398 420382 232634
rect 455826 232718 456062 232954
rect 456146 232718 456382 232954
rect 455826 232398 456062 232634
rect 456146 232398 456382 232634
rect 491826 232718 492062 232954
rect 492146 232718 492382 232954
rect 491826 232398 492062 232634
rect 492146 232398 492382 232634
rect 527826 232718 528062 232954
rect 528146 232718 528382 232954
rect 527826 232398 528062 232634
rect 528146 232398 528382 232634
rect 563826 232718 564062 232954
rect 564146 232718 564382 232954
rect 563826 232398 564062 232634
rect 564146 232398 564382 232634
rect 582326 232718 582562 232954
rect 582646 232718 582882 232954
rect 582326 232398 582562 232634
rect 582646 232398 582882 232634
rect -1974 228218 -1738 228454
rect -1654 228218 -1418 228454
rect -1974 227898 -1738 228134
rect -1654 227898 -1418 228134
rect 5826 228218 6062 228454
rect 6146 228218 6382 228454
rect 5826 227898 6062 228134
rect 6146 227898 6382 228134
rect 41826 228218 42062 228454
rect 42146 228218 42382 228454
rect 41826 227898 42062 228134
rect 42146 227898 42382 228134
rect 77826 228218 78062 228454
rect 78146 228218 78382 228454
rect 77826 227898 78062 228134
rect 78146 227898 78382 228134
rect 113826 228218 114062 228454
rect 114146 228218 114382 228454
rect 113826 227898 114062 228134
rect 114146 227898 114382 228134
rect 149826 228218 150062 228454
rect 150146 228218 150382 228454
rect 149826 227898 150062 228134
rect 150146 227898 150382 228134
rect 185826 228218 186062 228454
rect 186146 228218 186382 228454
rect 185826 227898 186062 228134
rect 186146 227898 186382 228134
rect 221826 228218 222062 228454
rect 222146 228218 222382 228454
rect 221826 227898 222062 228134
rect 222146 227898 222382 228134
rect 257826 228218 258062 228454
rect 258146 228218 258382 228454
rect 257826 227898 258062 228134
rect 258146 227898 258382 228134
rect 293826 228218 294062 228454
rect 294146 228218 294382 228454
rect 293826 227898 294062 228134
rect 294146 227898 294382 228134
rect 329826 228218 330062 228454
rect 330146 228218 330382 228454
rect 329826 227898 330062 228134
rect 330146 227898 330382 228134
rect 365826 228218 366062 228454
rect 366146 228218 366382 228454
rect 365826 227898 366062 228134
rect 366146 227898 366382 228134
rect 401826 228218 402062 228454
rect 402146 228218 402382 228454
rect 401826 227898 402062 228134
rect 402146 227898 402382 228134
rect 437826 228218 438062 228454
rect 438146 228218 438382 228454
rect 437826 227898 438062 228134
rect 438146 227898 438382 228134
rect 473826 228218 474062 228454
rect 474146 228218 474382 228454
rect 473826 227898 474062 228134
rect 474146 227898 474382 228134
rect 509826 228218 510062 228454
rect 510146 228218 510382 228454
rect 509826 227898 510062 228134
rect 510146 227898 510382 228134
rect 545826 228218 546062 228454
rect 546146 228218 546382 228454
rect 545826 227898 546062 228134
rect 546146 227898 546382 228134
rect 13198 196718 13434 196954
rect 13518 196718 13754 196954
rect 13198 196398 13434 196634
rect 13518 196398 13754 196634
rect 167826 196718 168062 196954
rect 168146 196718 168382 196954
rect 167826 196398 168062 196634
rect 168146 196398 168382 196634
rect 203826 196718 204062 196954
rect 204146 196718 204382 196954
rect 203826 196398 204062 196634
rect 204146 196398 204382 196634
rect 239826 196718 240062 196954
rect 240146 196718 240382 196954
rect 239826 196398 240062 196634
rect 240146 196398 240382 196634
rect 275826 196718 276062 196954
rect 276146 196718 276382 196954
rect 275826 196398 276062 196634
rect 276146 196398 276382 196634
rect 311826 196718 312062 196954
rect 312146 196718 312382 196954
rect 311826 196398 312062 196634
rect 312146 196398 312382 196634
rect 347826 196718 348062 196954
rect 348146 196718 348382 196954
rect 347826 196398 348062 196634
rect 348146 196398 348382 196634
rect 383826 196718 384062 196954
rect 384146 196718 384382 196954
rect 383826 196398 384062 196634
rect 384146 196398 384382 196634
rect 419826 196718 420062 196954
rect 420146 196718 420382 196954
rect 419826 196398 420062 196634
rect 420146 196398 420382 196634
rect 563826 196718 564062 196954
rect 564146 196718 564382 196954
rect 563826 196398 564062 196634
rect 564146 196398 564382 196634
rect 582326 196718 582562 196954
rect 582646 196718 582882 196954
rect 582326 196398 582562 196634
rect 582646 196398 582882 196634
rect -1974 192218 -1738 192454
rect -1654 192218 -1418 192454
rect -1974 191898 -1738 192134
rect -1654 191898 -1418 192134
rect 5826 192218 6062 192454
rect 6146 192218 6382 192454
rect 5826 191898 6062 192134
rect 6146 191898 6382 192134
rect 185826 192218 186062 192454
rect 186146 192218 186382 192454
rect 185826 191898 186062 192134
rect 186146 191898 186382 192134
rect 221826 192218 222062 192454
rect 222146 192218 222382 192454
rect 221826 191898 222062 192134
rect 222146 191898 222382 192134
rect 257826 192218 258062 192454
rect 258146 192218 258382 192454
rect 257826 191898 258062 192134
rect 258146 191898 258382 192134
rect 293826 192218 294062 192454
rect 294146 192218 294382 192454
rect 293826 191898 294062 192134
rect 294146 191898 294382 192134
rect 329826 192218 330062 192454
rect 330146 192218 330382 192454
rect 329826 191898 330062 192134
rect 330146 191898 330382 192134
rect 365826 192218 366062 192454
rect 366146 192218 366382 192454
rect 365826 191898 366062 192134
rect 366146 191898 366382 192134
rect 401826 192218 402062 192454
rect 402146 192218 402382 192454
rect 401826 191898 402062 192134
rect 402146 191898 402382 192134
rect 570350 192218 570586 192454
rect 570670 192218 570906 192454
rect 570350 191898 570586 192134
rect 570670 191898 570906 192134
rect 13198 160718 13434 160954
rect 13518 160718 13754 160954
rect 13198 160398 13434 160634
rect 13518 160398 13754 160634
rect 167826 160718 168062 160954
rect 168146 160718 168382 160954
rect 167826 160398 168062 160634
rect 168146 160398 168382 160634
rect 203826 160718 204062 160954
rect 204146 160718 204382 160954
rect 203826 160398 204062 160634
rect 204146 160398 204382 160634
rect 239826 160718 240062 160954
rect 240146 160718 240382 160954
rect 239826 160398 240062 160634
rect 240146 160398 240382 160634
rect 275826 160718 276062 160954
rect 276146 160718 276382 160954
rect 275826 160398 276062 160634
rect 276146 160398 276382 160634
rect 311826 160718 312062 160954
rect 312146 160718 312382 160954
rect 311826 160398 312062 160634
rect 312146 160398 312382 160634
rect 347826 160718 348062 160954
rect 348146 160718 348382 160954
rect 347826 160398 348062 160634
rect 348146 160398 348382 160634
rect 383826 160718 384062 160954
rect 384146 160718 384382 160954
rect 383826 160398 384062 160634
rect 384146 160398 384382 160634
rect 419826 160718 420062 160954
rect 420146 160718 420382 160954
rect 419826 160398 420062 160634
rect 420146 160398 420382 160634
rect 563826 160718 564062 160954
rect 564146 160718 564382 160954
rect 563826 160398 564062 160634
rect 564146 160398 564382 160634
rect 582326 160718 582562 160954
rect 582646 160718 582882 160954
rect 582326 160398 582562 160634
rect 582646 160398 582882 160634
rect -1974 156218 -1738 156454
rect -1654 156218 -1418 156454
rect -1974 155898 -1738 156134
rect -1654 155898 -1418 156134
rect 5826 156218 6062 156454
rect 6146 156218 6382 156454
rect 5826 155898 6062 156134
rect 6146 155898 6382 156134
rect 185826 156218 186062 156454
rect 186146 156218 186382 156454
rect 185826 155898 186062 156134
rect 186146 155898 186382 156134
rect 221826 156218 222062 156454
rect 222146 156218 222382 156454
rect 221826 155898 222062 156134
rect 222146 155898 222382 156134
rect 257826 156218 258062 156454
rect 258146 156218 258382 156454
rect 257826 155898 258062 156134
rect 258146 155898 258382 156134
rect 293826 156218 294062 156454
rect 294146 156218 294382 156454
rect 293826 155898 294062 156134
rect 294146 155898 294382 156134
rect 329826 156218 330062 156454
rect 330146 156218 330382 156454
rect 329826 155898 330062 156134
rect 330146 155898 330382 156134
rect 365826 156218 366062 156454
rect 366146 156218 366382 156454
rect 365826 155898 366062 156134
rect 366146 155898 366382 156134
rect 401826 156218 402062 156454
rect 402146 156218 402382 156454
rect 401826 155898 402062 156134
rect 402146 155898 402382 156134
rect 570350 156218 570586 156454
rect 570670 156218 570906 156454
rect 570350 155898 570586 156134
rect 570670 155898 570906 156134
rect 23826 124718 24062 124954
rect 24146 124718 24382 124954
rect 23826 124398 24062 124634
rect 24146 124398 24382 124634
rect 59826 124718 60062 124954
rect 60146 124718 60382 124954
rect 59826 124398 60062 124634
rect 60146 124398 60382 124634
rect 95826 124718 96062 124954
rect 96146 124718 96382 124954
rect 95826 124398 96062 124634
rect 96146 124398 96382 124634
rect 131826 124718 132062 124954
rect 132146 124718 132382 124954
rect 131826 124398 132062 124634
rect 132146 124398 132382 124634
rect 167826 124718 168062 124954
rect 168146 124718 168382 124954
rect 167826 124398 168062 124634
rect 168146 124398 168382 124634
rect 203826 124718 204062 124954
rect 204146 124718 204382 124954
rect 203826 124398 204062 124634
rect 204146 124398 204382 124634
rect 239826 124718 240062 124954
rect 240146 124718 240382 124954
rect 239826 124398 240062 124634
rect 240146 124398 240382 124634
rect 275826 124718 276062 124954
rect 276146 124718 276382 124954
rect 275826 124398 276062 124634
rect 276146 124398 276382 124634
rect 311826 124718 312062 124954
rect 312146 124718 312382 124954
rect 311826 124398 312062 124634
rect 312146 124398 312382 124634
rect 347826 124718 348062 124954
rect 348146 124718 348382 124954
rect 347826 124398 348062 124634
rect 348146 124398 348382 124634
rect 383826 124718 384062 124954
rect 384146 124718 384382 124954
rect 383826 124398 384062 124634
rect 384146 124398 384382 124634
rect 419826 124718 420062 124954
rect 420146 124718 420382 124954
rect 419826 124398 420062 124634
rect 420146 124398 420382 124634
rect 455826 124718 456062 124954
rect 456146 124718 456382 124954
rect 455826 124398 456062 124634
rect 456146 124398 456382 124634
rect 491826 124718 492062 124954
rect 492146 124718 492382 124954
rect 491826 124398 492062 124634
rect 492146 124398 492382 124634
rect 527826 124718 528062 124954
rect 528146 124718 528382 124954
rect 527826 124398 528062 124634
rect 528146 124398 528382 124634
rect 563826 124718 564062 124954
rect 564146 124718 564382 124954
rect 563826 124398 564062 124634
rect 564146 124398 564382 124634
rect 582326 124718 582562 124954
rect 582646 124718 582882 124954
rect 582326 124398 582562 124634
rect 582646 124398 582882 124634
rect -1974 120218 -1738 120454
rect -1654 120218 -1418 120454
rect -1974 119898 -1738 120134
rect -1654 119898 -1418 120134
rect 5826 120218 6062 120454
rect 6146 120218 6382 120454
rect 5826 119898 6062 120134
rect 6146 119898 6382 120134
rect 41826 120218 42062 120454
rect 42146 120218 42382 120454
rect 41826 119898 42062 120134
rect 42146 119898 42382 120134
rect 77826 120218 78062 120454
rect 78146 120218 78382 120454
rect 77826 119898 78062 120134
rect 78146 119898 78382 120134
rect 113826 120218 114062 120454
rect 114146 120218 114382 120454
rect 113826 119898 114062 120134
rect 114146 119898 114382 120134
rect 149826 120218 150062 120454
rect 150146 120218 150382 120454
rect 149826 119898 150062 120134
rect 150146 119898 150382 120134
rect 185826 120218 186062 120454
rect 186146 120218 186382 120454
rect 185826 119898 186062 120134
rect 186146 119898 186382 120134
rect 221826 120218 222062 120454
rect 222146 120218 222382 120454
rect 221826 119898 222062 120134
rect 222146 119898 222382 120134
rect 257826 120218 258062 120454
rect 258146 120218 258382 120454
rect 257826 119898 258062 120134
rect 258146 119898 258382 120134
rect 293826 120218 294062 120454
rect 294146 120218 294382 120454
rect 293826 119898 294062 120134
rect 294146 119898 294382 120134
rect 329826 120218 330062 120454
rect 330146 120218 330382 120454
rect 329826 119898 330062 120134
rect 330146 119898 330382 120134
rect 365826 120218 366062 120454
rect 366146 120218 366382 120454
rect 365826 119898 366062 120134
rect 366146 119898 366382 120134
rect 401826 120218 402062 120454
rect 402146 120218 402382 120454
rect 401826 119898 402062 120134
rect 402146 119898 402382 120134
rect 437826 120218 438062 120454
rect 438146 120218 438382 120454
rect 437826 119898 438062 120134
rect 438146 119898 438382 120134
rect 473826 120218 474062 120454
rect 474146 120218 474382 120454
rect 473826 119898 474062 120134
rect 474146 119898 474382 120134
rect 509826 120218 510062 120454
rect 510146 120218 510382 120454
rect 509826 119898 510062 120134
rect 510146 119898 510382 120134
rect 545826 120218 546062 120454
rect 546146 120218 546382 120454
rect 545826 119898 546062 120134
rect 546146 119898 546382 120134
rect 13198 88718 13434 88954
rect 13518 88718 13754 88954
rect 13198 88398 13434 88634
rect 13518 88398 13754 88634
rect 167826 88718 168062 88954
rect 168146 88718 168382 88954
rect 167826 88398 168062 88634
rect 168146 88398 168382 88634
rect 291590 88718 291826 88954
rect 291910 88718 292146 88954
rect 291590 88398 291826 88634
rect 291910 88398 292146 88634
rect 419826 88718 420062 88954
rect 420146 88718 420382 88954
rect 419826 88398 420062 88634
rect 420146 88398 420382 88634
rect 563826 88718 564062 88954
rect 564146 88718 564382 88954
rect 563826 88398 564062 88634
rect 564146 88398 564382 88634
rect 582326 88718 582562 88954
rect 582646 88718 582882 88954
rect 582326 88398 582562 88634
rect 582646 88398 582882 88634
rect -1974 84218 -1738 84454
rect -1654 84218 -1418 84454
rect -1974 83898 -1738 84134
rect -1654 83898 -1418 84134
rect 5826 84218 6062 84454
rect 6146 84218 6382 84454
rect 5826 83898 6062 84134
rect 6146 83898 6382 84134
rect 173094 84218 173330 84454
rect 173414 84218 173650 84454
rect 173094 83898 173330 84134
rect 173414 83898 173650 84134
rect 293826 84218 294062 84454
rect 294146 84218 294382 84454
rect 293826 83898 294062 84134
rect 294146 83898 294382 84134
rect 401826 84218 402062 84454
rect 402146 84218 402382 84454
rect 401826 83898 402062 84134
rect 402146 83898 402382 84134
rect 570350 84218 570586 84454
rect 570670 84218 570906 84454
rect 570350 83898 570586 84134
rect 570670 83898 570906 84134
rect 13198 52718 13434 52954
rect 13518 52718 13754 52954
rect 13198 52398 13434 52634
rect 13518 52398 13754 52634
rect 167826 52718 168062 52954
rect 168146 52718 168382 52954
rect 167826 52398 168062 52634
rect 168146 52398 168382 52634
rect 291590 52718 291826 52954
rect 291910 52718 292146 52954
rect 291590 52398 291826 52634
rect 291910 52398 292146 52634
rect 419826 52718 420062 52954
rect 420146 52718 420382 52954
rect 419826 52398 420062 52634
rect 420146 52398 420382 52634
rect 563826 52718 564062 52954
rect 564146 52718 564382 52954
rect 563826 52398 564062 52634
rect 564146 52398 564382 52634
rect 582326 52718 582562 52954
rect 582646 52718 582882 52954
rect 582326 52398 582562 52634
rect 582646 52398 582882 52634
rect -1974 48218 -1738 48454
rect -1654 48218 -1418 48454
rect -1974 47898 -1738 48134
rect -1654 47898 -1418 48134
rect 5826 48218 6062 48454
rect 6146 48218 6382 48454
rect 5826 47898 6062 48134
rect 6146 47898 6382 48134
rect 173094 48218 173330 48454
rect 173414 48218 173650 48454
rect 173094 47898 173330 48134
rect 173414 47898 173650 48134
rect 293826 48218 294062 48454
rect 294146 48218 294382 48454
rect 293826 47898 294062 48134
rect 294146 47898 294382 48134
rect 401826 48218 402062 48454
rect 402146 48218 402382 48454
rect 401826 47898 402062 48134
rect 402146 47898 402382 48134
rect 570350 48218 570586 48454
rect 570670 48218 570906 48454
rect 570350 47898 570586 48134
rect 570670 47898 570906 48134
rect 23826 16718 24062 16954
rect 24146 16718 24382 16954
rect 23826 16398 24062 16634
rect 24146 16398 24382 16634
rect 59826 16718 60062 16954
rect 60146 16718 60382 16954
rect 59826 16398 60062 16634
rect 60146 16398 60382 16634
rect 95826 16718 96062 16954
rect 96146 16718 96382 16954
rect 95826 16398 96062 16634
rect 96146 16398 96382 16634
rect 131826 16718 132062 16954
rect 132146 16718 132382 16954
rect 131826 16398 132062 16634
rect 132146 16398 132382 16634
rect 167826 16718 168062 16954
rect 168146 16718 168382 16954
rect 167826 16398 168062 16634
rect 168146 16398 168382 16634
rect 203826 16718 204062 16954
rect 204146 16718 204382 16954
rect 203826 16398 204062 16634
rect 204146 16398 204382 16634
rect 239826 16718 240062 16954
rect 240146 16718 240382 16954
rect 239826 16398 240062 16634
rect 240146 16398 240382 16634
rect 275826 16718 276062 16954
rect 276146 16718 276382 16954
rect 275826 16398 276062 16634
rect 276146 16398 276382 16634
rect 311826 16718 312062 16954
rect 312146 16718 312382 16954
rect 311826 16398 312062 16634
rect 312146 16398 312382 16634
rect 347826 16718 348062 16954
rect 348146 16718 348382 16954
rect 347826 16398 348062 16634
rect 348146 16398 348382 16634
rect 383826 16718 384062 16954
rect 384146 16718 384382 16954
rect 383826 16398 384062 16634
rect 384146 16398 384382 16634
rect 419826 16718 420062 16954
rect 420146 16718 420382 16954
rect 419826 16398 420062 16634
rect 420146 16398 420382 16634
rect 455826 16718 456062 16954
rect 456146 16718 456382 16954
rect 455826 16398 456062 16634
rect 456146 16398 456382 16634
rect 491826 16718 492062 16954
rect 492146 16718 492382 16954
rect 491826 16398 492062 16634
rect 492146 16398 492382 16634
rect 527826 16718 528062 16954
rect 528146 16718 528382 16954
rect 527826 16398 528062 16634
rect 528146 16398 528382 16634
rect 563826 16718 564062 16954
rect 564146 16718 564382 16954
rect 563826 16398 564062 16634
rect 564146 16398 564382 16634
rect 582326 16718 582562 16954
rect 582646 16718 582882 16954
rect 582326 16398 582562 16634
rect 582646 16398 582882 16634
rect -1974 12218 -1738 12454
rect -1654 12218 -1418 12454
rect -1974 11898 -1738 12134
rect -1654 11898 -1418 12134
rect 5826 12218 6062 12454
rect 6146 12218 6382 12454
rect 5826 11898 6062 12134
rect 6146 11898 6382 12134
rect 41826 12218 42062 12454
rect 42146 12218 42382 12454
rect 41826 11898 42062 12134
rect 42146 11898 42382 12134
rect 77826 12218 78062 12454
rect 78146 12218 78382 12454
rect 77826 11898 78062 12134
rect 78146 11898 78382 12134
rect 113826 12218 114062 12454
rect 114146 12218 114382 12454
rect 113826 11898 114062 12134
rect 114146 11898 114382 12134
rect 149826 12218 150062 12454
rect 150146 12218 150382 12454
rect 149826 11898 150062 12134
rect 150146 11898 150382 12134
rect 185826 12218 186062 12454
rect 186146 12218 186382 12454
rect 185826 11898 186062 12134
rect 186146 11898 186382 12134
rect 221826 12218 222062 12454
rect 222146 12218 222382 12454
rect 221826 11898 222062 12134
rect 222146 11898 222382 12134
rect 257826 12218 258062 12454
rect 258146 12218 258382 12454
rect 257826 11898 258062 12134
rect 258146 11898 258382 12134
rect 293826 12218 294062 12454
rect 294146 12218 294382 12454
rect 293826 11898 294062 12134
rect 294146 11898 294382 12134
rect 329826 12218 330062 12454
rect 330146 12218 330382 12454
rect 329826 11898 330062 12134
rect 330146 11898 330382 12134
rect 365826 12218 366062 12454
rect 366146 12218 366382 12454
rect 365826 11898 366062 12134
rect 366146 11898 366382 12134
rect 401826 12218 402062 12454
rect 402146 12218 402382 12454
rect 401826 11898 402062 12134
rect 402146 11898 402382 12134
rect 437826 12218 438062 12454
rect 438146 12218 438382 12454
rect 437826 11898 438062 12134
rect 438146 11898 438382 12134
rect 473826 12218 474062 12454
rect 474146 12218 474382 12454
rect 473826 11898 474062 12134
rect 474146 11898 474382 12134
rect 509826 12218 510062 12454
rect 510146 12218 510382 12454
rect 509826 11898 510062 12134
rect 510146 11898 510382 12134
rect 545826 12218 546062 12454
rect 546146 12218 546382 12454
rect 545826 11898 546062 12134
rect 546146 11898 546382 12134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 696218 585578 696454
rect 585662 696218 585898 696454
rect 585342 695898 585578 696134
rect 585662 695898 585898 696134
rect 585342 660218 585578 660454
rect 585662 660218 585898 660454
rect 585342 659898 585578 660134
rect 585662 659898 585898 660134
rect 585342 624218 585578 624454
rect 585662 624218 585898 624454
rect 585342 623898 585578 624134
rect 585662 623898 585898 624134
rect 585342 588218 585578 588454
rect 585662 588218 585898 588454
rect 585342 587898 585578 588134
rect 585662 587898 585898 588134
rect 585342 552218 585578 552454
rect 585662 552218 585898 552454
rect 585342 551898 585578 552134
rect 585662 551898 585898 552134
rect 585342 516218 585578 516454
rect 585662 516218 585898 516454
rect 585342 515898 585578 516134
rect 585662 515898 585898 516134
rect 585342 480218 585578 480454
rect 585662 480218 585898 480454
rect 585342 479898 585578 480134
rect 585662 479898 585898 480134
rect 585342 444218 585578 444454
rect 585662 444218 585898 444454
rect 585342 443898 585578 444134
rect 585662 443898 585898 444134
rect 585342 408218 585578 408454
rect 585662 408218 585898 408454
rect 585342 407898 585578 408134
rect 585662 407898 585898 408134
rect 585342 372218 585578 372454
rect 585662 372218 585898 372454
rect 585342 371898 585578 372134
rect 585662 371898 585898 372134
rect 585342 336218 585578 336454
rect 585662 336218 585898 336454
rect 585342 335898 585578 336134
rect 585662 335898 585898 336134
rect 585342 300218 585578 300454
rect 585662 300218 585898 300454
rect 585342 299898 585578 300134
rect 585662 299898 585898 300134
rect 585342 264218 585578 264454
rect 585662 264218 585898 264454
rect 585342 263898 585578 264134
rect 585662 263898 585898 264134
rect 585342 228218 585578 228454
rect 585662 228218 585898 228454
rect 585342 227898 585578 228134
rect 585662 227898 585898 228134
rect 585342 192218 585578 192454
rect 585662 192218 585898 192454
rect 585342 191898 585578 192134
rect 585662 191898 585898 192134
rect 585342 156218 585578 156454
rect 585662 156218 585898 156454
rect 585342 155898 585578 156134
rect 585662 155898 585898 156134
rect 585342 120218 585578 120454
rect 585662 120218 585898 120454
rect 585342 119898 585578 120134
rect 585662 119898 585898 120134
rect 585342 84218 585578 84454
rect 585662 84218 585898 84454
rect 585342 83898 585578 84134
rect 585662 83898 585898 84134
rect 585342 48218 585578 48454
rect 585662 48218 585898 48454
rect 585342 47898 585578 48134
rect 585662 47898 585898 48134
rect 585342 12218 585578 12454
rect 585662 12218 585898 12454
rect 585342 11898 585578 12134
rect 585662 11898 585898 12134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 700718 586538 700954
rect 586622 700718 586858 700954
rect 586302 700398 586538 700634
rect 586622 700398 586858 700634
rect 586302 664718 586538 664954
rect 586622 664718 586858 664954
rect 586302 664398 586538 664634
rect 586622 664398 586858 664634
rect 586302 628718 586538 628954
rect 586622 628718 586858 628954
rect 586302 628398 586538 628634
rect 586622 628398 586858 628634
rect 586302 592718 586538 592954
rect 586622 592718 586858 592954
rect 586302 592398 586538 592634
rect 586622 592398 586858 592634
rect 586302 556718 586538 556954
rect 586622 556718 586858 556954
rect 586302 556398 586538 556634
rect 586622 556398 586858 556634
rect 586302 520718 586538 520954
rect 586622 520718 586858 520954
rect 586302 520398 586538 520634
rect 586622 520398 586858 520634
rect 586302 484718 586538 484954
rect 586622 484718 586858 484954
rect 586302 484398 586538 484634
rect 586622 484398 586858 484634
rect 586302 448718 586538 448954
rect 586622 448718 586858 448954
rect 586302 448398 586538 448634
rect 586622 448398 586858 448634
rect 586302 412718 586538 412954
rect 586622 412718 586858 412954
rect 586302 412398 586538 412634
rect 586622 412398 586858 412634
rect 586302 376718 586538 376954
rect 586622 376718 586858 376954
rect 586302 376398 586538 376634
rect 586622 376398 586858 376634
rect 586302 340718 586538 340954
rect 586622 340718 586858 340954
rect 586302 340398 586538 340634
rect 586622 340398 586858 340634
rect 586302 304718 586538 304954
rect 586622 304718 586858 304954
rect 586302 304398 586538 304634
rect 586622 304398 586858 304634
rect 586302 268718 586538 268954
rect 586622 268718 586858 268954
rect 586302 268398 586538 268634
rect 586622 268398 586858 268634
rect 586302 232718 586538 232954
rect 586622 232718 586858 232954
rect 586302 232398 586538 232634
rect 586622 232398 586858 232634
rect 586302 196718 586538 196954
rect 586622 196718 586858 196954
rect 586302 196398 586538 196634
rect 586622 196398 586858 196634
rect 586302 160718 586538 160954
rect 586622 160718 586858 160954
rect 586302 160398 586538 160634
rect 586622 160398 586858 160634
rect 586302 124718 586538 124954
rect 586622 124718 586858 124954
rect 586302 124398 586538 124634
rect 586622 124398 586858 124634
rect 586302 88718 586538 88954
rect 586622 88718 586858 88954
rect 586302 88398 586538 88634
rect 586622 88398 586858 88634
rect 586302 52718 586538 52954
rect 586622 52718 586858 52954
rect 586302 52398 586538 52634
rect 586622 52398 586858 52634
rect 586302 16718 586538 16954
rect 586622 16718 586858 16954
rect 586302 16398 586538 16634
rect 586622 16398 586858 16634
rect 582326 -1542 582562 -1306
rect 582646 -1542 582882 -1306
rect 582326 -1862 582562 -1626
rect 582646 -1862 582882 -1626
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 582326 705798
rect 582562 705562 582646 705798
rect 582882 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 582326 705478
rect 582562 705242 582646 705478
rect 582882 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 700954 592650 700986
rect -8726 700718 -2934 700954
rect -2698 700718 -2614 700954
rect -2378 700718 582326 700954
rect 582562 700718 582646 700954
rect 582882 700718 586302 700954
rect 586538 700718 586622 700954
rect 586858 700718 592650 700954
rect -8726 700634 592650 700718
rect -8726 700398 -2934 700634
rect -2698 700398 -2614 700634
rect -2378 700398 582326 700634
rect 582562 700398 582646 700634
rect 582882 700398 586302 700634
rect 586538 700398 586622 700634
rect 586858 700398 592650 700634
rect -8726 700366 592650 700398
rect -8726 696454 592650 696486
rect -8726 696218 -1974 696454
rect -1738 696218 -1654 696454
rect -1418 696218 5826 696454
rect 6062 696218 6146 696454
rect 6382 696218 41826 696454
rect 42062 696218 42146 696454
rect 42382 696218 77826 696454
rect 78062 696218 78146 696454
rect 78382 696218 113826 696454
rect 114062 696218 114146 696454
rect 114382 696218 149826 696454
rect 150062 696218 150146 696454
rect 150382 696218 185826 696454
rect 186062 696218 186146 696454
rect 186382 696218 221826 696454
rect 222062 696218 222146 696454
rect 222382 696218 257826 696454
rect 258062 696218 258146 696454
rect 258382 696218 293826 696454
rect 294062 696218 294146 696454
rect 294382 696218 329826 696454
rect 330062 696218 330146 696454
rect 330382 696218 365826 696454
rect 366062 696218 366146 696454
rect 366382 696218 401826 696454
rect 402062 696218 402146 696454
rect 402382 696218 437826 696454
rect 438062 696218 438146 696454
rect 438382 696218 473826 696454
rect 474062 696218 474146 696454
rect 474382 696218 509826 696454
rect 510062 696218 510146 696454
rect 510382 696218 545826 696454
rect 546062 696218 546146 696454
rect 546382 696218 585342 696454
rect 585578 696218 585662 696454
rect 585898 696218 592650 696454
rect -8726 696134 592650 696218
rect -8726 695898 -1974 696134
rect -1738 695898 -1654 696134
rect -1418 695898 5826 696134
rect 6062 695898 6146 696134
rect 6382 695898 41826 696134
rect 42062 695898 42146 696134
rect 42382 695898 77826 696134
rect 78062 695898 78146 696134
rect 78382 695898 113826 696134
rect 114062 695898 114146 696134
rect 114382 695898 149826 696134
rect 150062 695898 150146 696134
rect 150382 695898 185826 696134
rect 186062 695898 186146 696134
rect 186382 695898 221826 696134
rect 222062 695898 222146 696134
rect 222382 695898 257826 696134
rect 258062 695898 258146 696134
rect 258382 695898 293826 696134
rect 294062 695898 294146 696134
rect 294382 695898 329826 696134
rect 330062 695898 330146 696134
rect 330382 695898 365826 696134
rect 366062 695898 366146 696134
rect 366382 695898 401826 696134
rect 402062 695898 402146 696134
rect 402382 695898 437826 696134
rect 438062 695898 438146 696134
rect 438382 695898 473826 696134
rect 474062 695898 474146 696134
rect 474382 695898 509826 696134
rect 510062 695898 510146 696134
rect 510382 695898 545826 696134
rect 546062 695898 546146 696134
rect 546382 695898 585342 696134
rect 585578 695898 585662 696134
rect 585898 695898 592650 696134
rect -8726 695866 592650 695898
rect -8726 664954 592650 664986
rect -8726 664718 -2934 664954
rect -2698 664718 -2614 664954
rect -2378 664718 13198 664954
rect 13434 664718 13518 664954
rect 13754 664718 167826 664954
rect 168062 664718 168146 664954
rect 168382 664718 291590 664954
rect 291826 664718 291910 664954
rect 292146 664718 419826 664954
rect 420062 664718 420146 664954
rect 420382 664718 563826 664954
rect 564062 664718 564146 664954
rect 564382 664718 582326 664954
rect 582562 664718 582646 664954
rect 582882 664718 586302 664954
rect 586538 664718 586622 664954
rect 586858 664718 592650 664954
rect -8726 664634 592650 664718
rect -8726 664398 -2934 664634
rect -2698 664398 -2614 664634
rect -2378 664398 13198 664634
rect 13434 664398 13518 664634
rect 13754 664398 167826 664634
rect 168062 664398 168146 664634
rect 168382 664398 291590 664634
rect 291826 664398 291910 664634
rect 292146 664398 419826 664634
rect 420062 664398 420146 664634
rect 420382 664398 563826 664634
rect 564062 664398 564146 664634
rect 564382 664398 582326 664634
rect 582562 664398 582646 664634
rect 582882 664398 586302 664634
rect 586538 664398 586622 664634
rect 586858 664398 592650 664634
rect -8726 664366 592650 664398
rect -8726 660454 592650 660486
rect -8726 660218 -1974 660454
rect -1738 660218 -1654 660454
rect -1418 660218 5826 660454
rect 6062 660218 6146 660454
rect 6382 660218 173094 660454
rect 173330 660218 173414 660454
rect 173650 660218 293826 660454
rect 294062 660218 294146 660454
rect 294382 660218 401826 660454
rect 402062 660218 402146 660454
rect 402382 660218 570350 660454
rect 570586 660218 570670 660454
rect 570906 660218 585342 660454
rect 585578 660218 585662 660454
rect 585898 660218 592650 660454
rect -8726 660134 592650 660218
rect -8726 659898 -1974 660134
rect -1738 659898 -1654 660134
rect -1418 659898 5826 660134
rect 6062 659898 6146 660134
rect 6382 659898 173094 660134
rect 173330 659898 173414 660134
rect 173650 659898 293826 660134
rect 294062 659898 294146 660134
rect 294382 659898 401826 660134
rect 402062 659898 402146 660134
rect 402382 659898 570350 660134
rect 570586 659898 570670 660134
rect 570906 659898 585342 660134
rect 585578 659898 585662 660134
rect 585898 659898 592650 660134
rect -8726 659866 592650 659898
rect -8726 628954 592650 628986
rect -8726 628718 -2934 628954
rect -2698 628718 -2614 628954
rect -2378 628718 13198 628954
rect 13434 628718 13518 628954
rect 13754 628718 167826 628954
rect 168062 628718 168146 628954
rect 168382 628718 291590 628954
rect 291826 628718 291910 628954
rect 292146 628718 419826 628954
rect 420062 628718 420146 628954
rect 420382 628718 563826 628954
rect 564062 628718 564146 628954
rect 564382 628718 582326 628954
rect 582562 628718 582646 628954
rect 582882 628718 586302 628954
rect 586538 628718 586622 628954
rect 586858 628718 592650 628954
rect -8726 628634 592650 628718
rect -8726 628398 -2934 628634
rect -2698 628398 -2614 628634
rect -2378 628398 13198 628634
rect 13434 628398 13518 628634
rect 13754 628398 167826 628634
rect 168062 628398 168146 628634
rect 168382 628398 291590 628634
rect 291826 628398 291910 628634
rect 292146 628398 419826 628634
rect 420062 628398 420146 628634
rect 420382 628398 563826 628634
rect 564062 628398 564146 628634
rect 564382 628398 582326 628634
rect 582562 628398 582646 628634
rect 582882 628398 586302 628634
rect 586538 628398 586622 628634
rect 586858 628398 592650 628634
rect -8726 628366 592650 628398
rect -8726 624454 592650 624486
rect -8726 624218 -1974 624454
rect -1738 624218 -1654 624454
rect -1418 624218 5826 624454
rect 6062 624218 6146 624454
rect 6382 624218 173094 624454
rect 173330 624218 173414 624454
rect 173650 624218 293826 624454
rect 294062 624218 294146 624454
rect 294382 624218 401826 624454
rect 402062 624218 402146 624454
rect 402382 624218 570350 624454
rect 570586 624218 570670 624454
rect 570906 624218 585342 624454
rect 585578 624218 585662 624454
rect 585898 624218 592650 624454
rect -8726 624134 592650 624218
rect -8726 623898 -1974 624134
rect -1738 623898 -1654 624134
rect -1418 623898 5826 624134
rect 6062 623898 6146 624134
rect 6382 623898 173094 624134
rect 173330 623898 173414 624134
rect 173650 623898 293826 624134
rect 294062 623898 294146 624134
rect 294382 623898 401826 624134
rect 402062 623898 402146 624134
rect 402382 623898 570350 624134
rect 570586 623898 570670 624134
rect 570906 623898 585342 624134
rect 585578 623898 585662 624134
rect 585898 623898 592650 624134
rect -8726 623866 592650 623898
rect -8726 592954 592650 592986
rect -8726 592718 -2934 592954
rect -2698 592718 -2614 592954
rect -2378 592718 23826 592954
rect 24062 592718 24146 592954
rect 24382 592718 59826 592954
rect 60062 592718 60146 592954
rect 60382 592718 95826 592954
rect 96062 592718 96146 592954
rect 96382 592718 131826 592954
rect 132062 592718 132146 592954
rect 132382 592718 167826 592954
rect 168062 592718 168146 592954
rect 168382 592718 291590 592954
rect 291826 592718 291910 592954
rect 292146 592718 419826 592954
rect 420062 592718 420146 592954
rect 420382 592718 455826 592954
rect 456062 592718 456146 592954
rect 456382 592718 491826 592954
rect 492062 592718 492146 592954
rect 492382 592718 527826 592954
rect 528062 592718 528146 592954
rect 528382 592718 563826 592954
rect 564062 592718 564146 592954
rect 564382 592718 582326 592954
rect 582562 592718 582646 592954
rect 582882 592718 586302 592954
rect 586538 592718 586622 592954
rect 586858 592718 592650 592954
rect -8726 592634 592650 592718
rect -8726 592398 -2934 592634
rect -2698 592398 -2614 592634
rect -2378 592398 23826 592634
rect 24062 592398 24146 592634
rect 24382 592398 59826 592634
rect 60062 592398 60146 592634
rect 60382 592398 95826 592634
rect 96062 592398 96146 592634
rect 96382 592398 131826 592634
rect 132062 592398 132146 592634
rect 132382 592398 167826 592634
rect 168062 592398 168146 592634
rect 168382 592398 291590 592634
rect 291826 592398 291910 592634
rect 292146 592398 419826 592634
rect 420062 592398 420146 592634
rect 420382 592398 455826 592634
rect 456062 592398 456146 592634
rect 456382 592398 491826 592634
rect 492062 592398 492146 592634
rect 492382 592398 527826 592634
rect 528062 592398 528146 592634
rect 528382 592398 563826 592634
rect 564062 592398 564146 592634
rect 564382 592398 582326 592634
rect 582562 592398 582646 592634
rect 582882 592398 586302 592634
rect 586538 592398 586622 592634
rect 586858 592398 592650 592634
rect -8726 592366 592650 592398
rect -8726 588454 592650 588486
rect -8726 588218 -1974 588454
rect -1738 588218 -1654 588454
rect -1418 588218 5826 588454
rect 6062 588218 6146 588454
rect 6382 588218 41826 588454
rect 42062 588218 42146 588454
rect 42382 588218 77826 588454
rect 78062 588218 78146 588454
rect 78382 588218 113826 588454
rect 114062 588218 114146 588454
rect 114382 588218 149826 588454
rect 150062 588218 150146 588454
rect 150382 588218 185826 588454
rect 186062 588218 186146 588454
rect 186382 588218 221826 588454
rect 222062 588218 222146 588454
rect 222382 588218 257826 588454
rect 258062 588218 258146 588454
rect 258382 588218 293826 588454
rect 294062 588218 294146 588454
rect 294382 588218 329826 588454
rect 330062 588218 330146 588454
rect 330382 588218 365826 588454
rect 366062 588218 366146 588454
rect 366382 588218 401826 588454
rect 402062 588218 402146 588454
rect 402382 588218 437826 588454
rect 438062 588218 438146 588454
rect 438382 588218 473826 588454
rect 474062 588218 474146 588454
rect 474382 588218 509826 588454
rect 510062 588218 510146 588454
rect 510382 588218 545826 588454
rect 546062 588218 546146 588454
rect 546382 588218 585342 588454
rect 585578 588218 585662 588454
rect 585898 588218 592650 588454
rect -8726 588134 592650 588218
rect -8726 587898 -1974 588134
rect -1738 587898 -1654 588134
rect -1418 587898 5826 588134
rect 6062 587898 6146 588134
rect 6382 587898 41826 588134
rect 42062 587898 42146 588134
rect 42382 587898 77826 588134
rect 78062 587898 78146 588134
rect 78382 587898 113826 588134
rect 114062 587898 114146 588134
rect 114382 587898 149826 588134
rect 150062 587898 150146 588134
rect 150382 587898 185826 588134
rect 186062 587898 186146 588134
rect 186382 587898 221826 588134
rect 222062 587898 222146 588134
rect 222382 587898 257826 588134
rect 258062 587898 258146 588134
rect 258382 587898 293826 588134
rect 294062 587898 294146 588134
rect 294382 587898 329826 588134
rect 330062 587898 330146 588134
rect 330382 587898 365826 588134
rect 366062 587898 366146 588134
rect 366382 587898 401826 588134
rect 402062 587898 402146 588134
rect 402382 587898 437826 588134
rect 438062 587898 438146 588134
rect 438382 587898 473826 588134
rect 474062 587898 474146 588134
rect 474382 587898 509826 588134
rect 510062 587898 510146 588134
rect 510382 587898 545826 588134
rect 546062 587898 546146 588134
rect 546382 587898 585342 588134
rect 585578 587898 585662 588134
rect 585898 587898 592650 588134
rect -8726 587866 592650 587898
rect -8726 556954 592650 556986
rect -8726 556718 -2934 556954
rect -2698 556718 -2614 556954
rect -2378 556718 13198 556954
rect 13434 556718 13518 556954
rect 13754 556718 167826 556954
rect 168062 556718 168146 556954
rect 168382 556718 203826 556954
rect 204062 556718 204146 556954
rect 204382 556718 239826 556954
rect 240062 556718 240146 556954
rect 240382 556718 275826 556954
rect 276062 556718 276146 556954
rect 276382 556718 311826 556954
rect 312062 556718 312146 556954
rect 312382 556718 347826 556954
rect 348062 556718 348146 556954
rect 348382 556718 383826 556954
rect 384062 556718 384146 556954
rect 384382 556718 419826 556954
rect 420062 556718 420146 556954
rect 420382 556718 563826 556954
rect 564062 556718 564146 556954
rect 564382 556718 582326 556954
rect 582562 556718 582646 556954
rect 582882 556718 586302 556954
rect 586538 556718 586622 556954
rect 586858 556718 592650 556954
rect -8726 556634 592650 556718
rect -8726 556398 -2934 556634
rect -2698 556398 -2614 556634
rect -2378 556398 13198 556634
rect 13434 556398 13518 556634
rect 13754 556398 167826 556634
rect 168062 556398 168146 556634
rect 168382 556398 203826 556634
rect 204062 556398 204146 556634
rect 204382 556398 239826 556634
rect 240062 556398 240146 556634
rect 240382 556398 275826 556634
rect 276062 556398 276146 556634
rect 276382 556398 311826 556634
rect 312062 556398 312146 556634
rect 312382 556398 347826 556634
rect 348062 556398 348146 556634
rect 348382 556398 383826 556634
rect 384062 556398 384146 556634
rect 384382 556398 419826 556634
rect 420062 556398 420146 556634
rect 420382 556398 563826 556634
rect 564062 556398 564146 556634
rect 564382 556398 582326 556634
rect 582562 556398 582646 556634
rect 582882 556398 586302 556634
rect 586538 556398 586622 556634
rect 586858 556398 592650 556634
rect -8726 556366 592650 556398
rect -8726 552454 592650 552486
rect -8726 552218 -1974 552454
rect -1738 552218 -1654 552454
rect -1418 552218 5826 552454
rect 6062 552218 6146 552454
rect 6382 552218 185826 552454
rect 186062 552218 186146 552454
rect 186382 552218 221826 552454
rect 222062 552218 222146 552454
rect 222382 552218 257826 552454
rect 258062 552218 258146 552454
rect 258382 552218 293826 552454
rect 294062 552218 294146 552454
rect 294382 552218 329826 552454
rect 330062 552218 330146 552454
rect 330382 552218 365826 552454
rect 366062 552218 366146 552454
rect 366382 552218 401826 552454
rect 402062 552218 402146 552454
rect 402382 552218 570350 552454
rect 570586 552218 570670 552454
rect 570906 552218 585342 552454
rect 585578 552218 585662 552454
rect 585898 552218 592650 552454
rect -8726 552134 592650 552218
rect -8726 551898 -1974 552134
rect -1738 551898 -1654 552134
rect -1418 551898 5826 552134
rect 6062 551898 6146 552134
rect 6382 551898 185826 552134
rect 186062 551898 186146 552134
rect 186382 551898 221826 552134
rect 222062 551898 222146 552134
rect 222382 551898 257826 552134
rect 258062 551898 258146 552134
rect 258382 551898 293826 552134
rect 294062 551898 294146 552134
rect 294382 551898 329826 552134
rect 330062 551898 330146 552134
rect 330382 551898 365826 552134
rect 366062 551898 366146 552134
rect 366382 551898 401826 552134
rect 402062 551898 402146 552134
rect 402382 551898 570350 552134
rect 570586 551898 570670 552134
rect 570906 551898 585342 552134
rect 585578 551898 585662 552134
rect 585898 551898 592650 552134
rect -8726 551866 592650 551898
rect -8726 520954 592650 520986
rect -8726 520718 -2934 520954
rect -2698 520718 -2614 520954
rect -2378 520718 13198 520954
rect 13434 520718 13518 520954
rect 13754 520718 167826 520954
rect 168062 520718 168146 520954
rect 168382 520718 203826 520954
rect 204062 520718 204146 520954
rect 204382 520718 239826 520954
rect 240062 520718 240146 520954
rect 240382 520718 275826 520954
rect 276062 520718 276146 520954
rect 276382 520718 311826 520954
rect 312062 520718 312146 520954
rect 312382 520718 347826 520954
rect 348062 520718 348146 520954
rect 348382 520718 383826 520954
rect 384062 520718 384146 520954
rect 384382 520718 419826 520954
rect 420062 520718 420146 520954
rect 420382 520718 563826 520954
rect 564062 520718 564146 520954
rect 564382 520718 582326 520954
rect 582562 520718 582646 520954
rect 582882 520718 586302 520954
rect 586538 520718 586622 520954
rect 586858 520718 592650 520954
rect -8726 520634 592650 520718
rect -8726 520398 -2934 520634
rect -2698 520398 -2614 520634
rect -2378 520398 13198 520634
rect 13434 520398 13518 520634
rect 13754 520398 167826 520634
rect 168062 520398 168146 520634
rect 168382 520398 203826 520634
rect 204062 520398 204146 520634
rect 204382 520398 239826 520634
rect 240062 520398 240146 520634
rect 240382 520398 275826 520634
rect 276062 520398 276146 520634
rect 276382 520398 311826 520634
rect 312062 520398 312146 520634
rect 312382 520398 347826 520634
rect 348062 520398 348146 520634
rect 348382 520398 383826 520634
rect 384062 520398 384146 520634
rect 384382 520398 419826 520634
rect 420062 520398 420146 520634
rect 420382 520398 563826 520634
rect 564062 520398 564146 520634
rect 564382 520398 582326 520634
rect 582562 520398 582646 520634
rect 582882 520398 586302 520634
rect 586538 520398 586622 520634
rect 586858 520398 592650 520634
rect -8726 520366 592650 520398
rect -8726 516454 592650 516486
rect -8726 516218 -1974 516454
rect -1738 516218 -1654 516454
rect -1418 516218 5826 516454
rect 6062 516218 6146 516454
rect 6382 516218 185826 516454
rect 186062 516218 186146 516454
rect 186382 516218 221826 516454
rect 222062 516218 222146 516454
rect 222382 516218 257826 516454
rect 258062 516218 258146 516454
rect 258382 516218 293826 516454
rect 294062 516218 294146 516454
rect 294382 516218 329826 516454
rect 330062 516218 330146 516454
rect 330382 516218 365826 516454
rect 366062 516218 366146 516454
rect 366382 516218 401826 516454
rect 402062 516218 402146 516454
rect 402382 516218 570350 516454
rect 570586 516218 570670 516454
rect 570906 516218 585342 516454
rect 585578 516218 585662 516454
rect 585898 516218 592650 516454
rect -8726 516134 592650 516218
rect -8726 515898 -1974 516134
rect -1738 515898 -1654 516134
rect -1418 515898 5826 516134
rect 6062 515898 6146 516134
rect 6382 515898 185826 516134
rect 186062 515898 186146 516134
rect 186382 515898 221826 516134
rect 222062 515898 222146 516134
rect 222382 515898 257826 516134
rect 258062 515898 258146 516134
rect 258382 515898 293826 516134
rect 294062 515898 294146 516134
rect 294382 515898 329826 516134
rect 330062 515898 330146 516134
rect 330382 515898 365826 516134
rect 366062 515898 366146 516134
rect 366382 515898 401826 516134
rect 402062 515898 402146 516134
rect 402382 515898 570350 516134
rect 570586 515898 570670 516134
rect 570906 515898 585342 516134
rect 585578 515898 585662 516134
rect 585898 515898 592650 516134
rect -8726 515866 592650 515898
rect -8726 484954 592650 484986
rect -8726 484718 -2934 484954
rect -2698 484718 -2614 484954
rect -2378 484718 23826 484954
rect 24062 484718 24146 484954
rect 24382 484718 59826 484954
rect 60062 484718 60146 484954
rect 60382 484718 95826 484954
rect 96062 484718 96146 484954
rect 96382 484718 131826 484954
rect 132062 484718 132146 484954
rect 132382 484718 167826 484954
rect 168062 484718 168146 484954
rect 168382 484718 203826 484954
rect 204062 484718 204146 484954
rect 204382 484718 239826 484954
rect 240062 484718 240146 484954
rect 240382 484718 275826 484954
rect 276062 484718 276146 484954
rect 276382 484718 311826 484954
rect 312062 484718 312146 484954
rect 312382 484718 347826 484954
rect 348062 484718 348146 484954
rect 348382 484718 383826 484954
rect 384062 484718 384146 484954
rect 384382 484718 419826 484954
rect 420062 484718 420146 484954
rect 420382 484718 455826 484954
rect 456062 484718 456146 484954
rect 456382 484718 491826 484954
rect 492062 484718 492146 484954
rect 492382 484718 527826 484954
rect 528062 484718 528146 484954
rect 528382 484718 563826 484954
rect 564062 484718 564146 484954
rect 564382 484718 582326 484954
rect 582562 484718 582646 484954
rect 582882 484718 586302 484954
rect 586538 484718 586622 484954
rect 586858 484718 592650 484954
rect -8726 484634 592650 484718
rect -8726 484398 -2934 484634
rect -2698 484398 -2614 484634
rect -2378 484398 23826 484634
rect 24062 484398 24146 484634
rect 24382 484398 59826 484634
rect 60062 484398 60146 484634
rect 60382 484398 95826 484634
rect 96062 484398 96146 484634
rect 96382 484398 131826 484634
rect 132062 484398 132146 484634
rect 132382 484398 167826 484634
rect 168062 484398 168146 484634
rect 168382 484398 203826 484634
rect 204062 484398 204146 484634
rect 204382 484398 239826 484634
rect 240062 484398 240146 484634
rect 240382 484398 275826 484634
rect 276062 484398 276146 484634
rect 276382 484398 311826 484634
rect 312062 484398 312146 484634
rect 312382 484398 347826 484634
rect 348062 484398 348146 484634
rect 348382 484398 383826 484634
rect 384062 484398 384146 484634
rect 384382 484398 419826 484634
rect 420062 484398 420146 484634
rect 420382 484398 455826 484634
rect 456062 484398 456146 484634
rect 456382 484398 491826 484634
rect 492062 484398 492146 484634
rect 492382 484398 527826 484634
rect 528062 484398 528146 484634
rect 528382 484398 563826 484634
rect 564062 484398 564146 484634
rect 564382 484398 582326 484634
rect 582562 484398 582646 484634
rect 582882 484398 586302 484634
rect 586538 484398 586622 484634
rect 586858 484398 592650 484634
rect -8726 484366 592650 484398
rect -8726 480454 592650 480486
rect -8726 480218 -1974 480454
rect -1738 480218 -1654 480454
rect -1418 480218 5826 480454
rect 6062 480218 6146 480454
rect 6382 480218 41826 480454
rect 42062 480218 42146 480454
rect 42382 480218 77826 480454
rect 78062 480218 78146 480454
rect 78382 480218 113826 480454
rect 114062 480218 114146 480454
rect 114382 480218 149826 480454
rect 150062 480218 150146 480454
rect 150382 480218 185826 480454
rect 186062 480218 186146 480454
rect 186382 480218 221826 480454
rect 222062 480218 222146 480454
rect 222382 480218 257826 480454
rect 258062 480218 258146 480454
rect 258382 480218 293826 480454
rect 294062 480218 294146 480454
rect 294382 480218 329826 480454
rect 330062 480218 330146 480454
rect 330382 480218 365826 480454
rect 366062 480218 366146 480454
rect 366382 480218 401826 480454
rect 402062 480218 402146 480454
rect 402382 480218 437826 480454
rect 438062 480218 438146 480454
rect 438382 480218 473826 480454
rect 474062 480218 474146 480454
rect 474382 480218 509826 480454
rect 510062 480218 510146 480454
rect 510382 480218 545826 480454
rect 546062 480218 546146 480454
rect 546382 480218 585342 480454
rect 585578 480218 585662 480454
rect 585898 480218 592650 480454
rect -8726 480134 592650 480218
rect -8726 479898 -1974 480134
rect -1738 479898 -1654 480134
rect -1418 479898 5826 480134
rect 6062 479898 6146 480134
rect 6382 479898 41826 480134
rect 42062 479898 42146 480134
rect 42382 479898 77826 480134
rect 78062 479898 78146 480134
rect 78382 479898 113826 480134
rect 114062 479898 114146 480134
rect 114382 479898 149826 480134
rect 150062 479898 150146 480134
rect 150382 479898 185826 480134
rect 186062 479898 186146 480134
rect 186382 479898 221826 480134
rect 222062 479898 222146 480134
rect 222382 479898 257826 480134
rect 258062 479898 258146 480134
rect 258382 479898 293826 480134
rect 294062 479898 294146 480134
rect 294382 479898 329826 480134
rect 330062 479898 330146 480134
rect 330382 479898 365826 480134
rect 366062 479898 366146 480134
rect 366382 479898 401826 480134
rect 402062 479898 402146 480134
rect 402382 479898 437826 480134
rect 438062 479898 438146 480134
rect 438382 479898 473826 480134
rect 474062 479898 474146 480134
rect 474382 479898 509826 480134
rect 510062 479898 510146 480134
rect 510382 479898 545826 480134
rect 546062 479898 546146 480134
rect 546382 479898 585342 480134
rect 585578 479898 585662 480134
rect 585898 479898 592650 480134
rect -8726 479866 592650 479898
rect -8726 448954 592650 448986
rect -8726 448718 -2934 448954
rect -2698 448718 -2614 448954
rect -2378 448718 13198 448954
rect 13434 448718 13518 448954
rect 13754 448718 167826 448954
rect 168062 448718 168146 448954
rect 168382 448718 203826 448954
rect 204062 448718 204146 448954
rect 204382 448718 239826 448954
rect 240062 448718 240146 448954
rect 240382 448718 275826 448954
rect 276062 448718 276146 448954
rect 276382 448718 311826 448954
rect 312062 448718 312146 448954
rect 312382 448718 347826 448954
rect 348062 448718 348146 448954
rect 348382 448718 383826 448954
rect 384062 448718 384146 448954
rect 384382 448718 419826 448954
rect 420062 448718 420146 448954
rect 420382 448718 563826 448954
rect 564062 448718 564146 448954
rect 564382 448718 582326 448954
rect 582562 448718 582646 448954
rect 582882 448718 586302 448954
rect 586538 448718 586622 448954
rect 586858 448718 592650 448954
rect -8726 448634 592650 448718
rect -8726 448398 -2934 448634
rect -2698 448398 -2614 448634
rect -2378 448398 13198 448634
rect 13434 448398 13518 448634
rect 13754 448398 167826 448634
rect 168062 448398 168146 448634
rect 168382 448398 203826 448634
rect 204062 448398 204146 448634
rect 204382 448398 239826 448634
rect 240062 448398 240146 448634
rect 240382 448398 275826 448634
rect 276062 448398 276146 448634
rect 276382 448398 311826 448634
rect 312062 448398 312146 448634
rect 312382 448398 347826 448634
rect 348062 448398 348146 448634
rect 348382 448398 383826 448634
rect 384062 448398 384146 448634
rect 384382 448398 419826 448634
rect 420062 448398 420146 448634
rect 420382 448398 563826 448634
rect 564062 448398 564146 448634
rect 564382 448398 582326 448634
rect 582562 448398 582646 448634
rect 582882 448398 586302 448634
rect 586538 448398 586622 448634
rect 586858 448398 592650 448634
rect -8726 448366 592650 448398
rect -8726 444454 592650 444486
rect -8726 444218 -1974 444454
rect -1738 444218 -1654 444454
rect -1418 444218 5826 444454
rect 6062 444218 6146 444454
rect 6382 444218 185826 444454
rect 186062 444218 186146 444454
rect 186382 444218 221826 444454
rect 222062 444218 222146 444454
rect 222382 444218 257826 444454
rect 258062 444218 258146 444454
rect 258382 444218 293826 444454
rect 294062 444218 294146 444454
rect 294382 444218 329826 444454
rect 330062 444218 330146 444454
rect 330382 444218 365826 444454
rect 366062 444218 366146 444454
rect 366382 444218 401826 444454
rect 402062 444218 402146 444454
rect 402382 444218 570350 444454
rect 570586 444218 570670 444454
rect 570906 444218 585342 444454
rect 585578 444218 585662 444454
rect 585898 444218 592650 444454
rect -8726 444134 592650 444218
rect -8726 443898 -1974 444134
rect -1738 443898 -1654 444134
rect -1418 443898 5826 444134
rect 6062 443898 6146 444134
rect 6382 443898 185826 444134
rect 186062 443898 186146 444134
rect 186382 443898 221826 444134
rect 222062 443898 222146 444134
rect 222382 443898 257826 444134
rect 258062 443898 258146 444134
rect 258382 443898 293826 444134
rect 294062 443898 294146 444134
rect 294382 443898 329826 444134
rect 330062 443898 330146 444134
rect 330382 443898 365826 444134
rect 366062 443898 366146 444134
rect 366382 443898 401826 444134
rect 402062 443898 402146 444134
rect 402382 443898 570350 444134
rect 570586 443898 570670 444134
rect 570906 443898 585342 444134
rect 585578 443898 585662 444134
rect 585898 443898 592650 444134
rect -8726 443866 592650 443898
rect -8726 412954 592650 412986
rect -8726 412718 -2934 412954
rect -2698 412718 -2614 412954
rect -2378 412718 13198 412954
rect 13434 412718 13518 412954
rect 13754 412718 167826 412954
rect 168062 412718 168146 412954
rect 168382 412718 203826 412954
rect 204062 412718 204146 412954
rect 204382 412718 239826 412954
rect 240062 412718 240146 412954
rect 240382 412718 275826 412954
rect 276062 412718 276146 412954
rect 276382 412718 311826 412954
rect 312062 412718 312146 412954
rect 312382 412718 347826 412954
rect 348062 412718 348146 412954
rect 348382 412718 383826 412954
rect 384062 412718 384146 412954
rect 384382 412718 419826 412954
rect 420062 412718 420146 412954
rect 420382 412718 563826 412954
rect 564062 412718 564146 412954
rect 564382 412718 582326 412954
rect 582562 412718 582646 412954
rect 582882 412718 586302 412954
rect 586538 412718 586622 412954
rect 586858 412718 592650 412954
rect -8726 412634 592650 412718
rect -8726 412398 -2934 412634
rect -2698 412398 -2614 412634
rect -2378 412398 13198 412634
rect 13434 412398 13518 412634
rect 13754 412398 167826 412634
rect 168062 412398 168146 412634
rect 168382 412398 203826 412634
rect 204062 412398 204146 412634
rect 204382 412398 239826 412634
rect 240062 412398 240146 412634
rect 240382 412398 275826 412634
rect 276062 412398 276146 412634
rect 276382 412398 311826 412634
rect 312062 412398 312146 412634
rect 312382 412398 347826 412634
rect 348062 412398 348146 412634
rect 348382 412398 383826 412634
rect 384062 412398 384146 412634
rect 384382 412398 419826 412634
rect 420062 412398 420146 412634
rect 420382 412398 563826 412634
rect 564062 412398 564146 412634
rect 564382 412398 582326 412634
rect 582562 412398 582646 412634
rect 582882 412398 586302 412634
rect 586538 412398 586622 412634
rect 586858 412398 592650 412634
rect -8726 412366 592650 412398
rect -8726 408454 592650 408486
rect -8726 408218 -1974 408454
rect -1738 408218 -1654 408454
rect -1418 408218 5826 408454
rect 6062 408218 6146 408454
rect 6382 408218 185826 408454
rect 186062 408218 186146 408454
rect 186382 408218 221826 408454
rect 222062 408218 222146 408454
rect 222382 408218 257826 408454
rect 258062 408218 258146 408454
rect 258382 408218 293826 408454
rect 294062 408218 294146 408454
rect 294382 408218 329826 408454
rect 330062 408218 330146 408454
rect 330382 408218 365826 408454
rect 366062 408218 366146 408454
rect 366382 408218 401826 408454
rect 402062 408218 402146 408454
rect 402382 408218 570350 408454
rect 570586 408218 570670 408454
rect 570906 408218 585342 408454
rect 585578 408218 585662 408454
rect 585898 408218 592650 408454
rect -8726 408134 592650 408218
rect -8726 407898 -1974 408134
rect -1738 407898 -1654 408134
rect -1418 407898 5826 408134
rect 6062 407898 6146 408134
rect 6382 407898 185826 408134
rect 186062 407898 186146 408134
rect 186382 407898 221826 408134
rect 222062 407898 222146 408134
rect 222382 407898 257826 408134
rect 258062 407898 258146 408134
rect 258382 407898 293826 408134
rect 294062 407898 294146 408134
rect 294382 407898 329826 408134
rect 330062 407898 330146 408134
rect 330382 407898 365826 408134
rect 366062 407898 366146 408134
rect 366382 407898 401826 408134
rect 402062 407898 402146 408134
rect 402382 407898 570350 408134
rect 570586 407898 570670 408134
rect 570906 407898 585342 408134
rect 585578 407898 585662 408134
rect 585898 407898 592650 408134
rect -8726 407866 592650 407898
rect -8726 376954 592650 376986
rect -8726 376718 -2934 376954
rect -2698 376718 -2614 376954
rect -2378 376718 13198 376954
rect 13434 376718 13518 376954
rect 13754 376718 167826 376954
rect 168062 376718 168146 376954
rect 168382 376718 203826 376954
rect 204062 376718 204146 376954
rect 204382 376718 239826 376954
rect 240062 376718 240146 376954
rect 240382 376718 275826 376954
rect 276062 376718 276146 376954
rect 276382 376718 311826 376954
rect 312062 376718 312146 376954
rect 312382 376718 347826 376954
rect 348062 376718 348146 376954
rect 348382 376718 383826 376954
rect 384062 376718 384146 376954
rect 384382 376718 419826 376954
rect 420062 376718 420146 376954
rect 420382 376718 563826 376954
rect 564062 376718 564146 376954
rect 564382 376718 582326 376954
rect 582562 376718 582646 376954
rect 582882 376718 586302 376954
rect 586538 376718 586622 376954
rect 586858 376718 592650 376954
rect -8726 376634 592650 376718
rect -8726 376398 -2934 376634
rect -2698 376398 -2614 376634
rect -2378 376398 13198 376634
rect 13434 376398 13518 376634
rect 13754 376398 167826 376634
rect 168062 376398 168146 376634
rect 168382 376398 203826 376634
rect 204062 376398 204146 376634
rect 204382 376398 239826 376634
rect 240062 376398 240146 376634
rect 240382 376398 275826 376634
rect 276062 376398 276146 376634
rect 276382 376398 311826 376634
rect 312062 376398 312146 376634
rect 312382 376398 347826 376634
rect 348062 376398 348146 376634
rect 348382 376398 383826 376634
rect 384062 376398 384146 376634
rect 384382 376398 419826 376634
rect 420062 376398 420146 376634
rect 420382 376398 563826 376634
rect 564062 376398 564146 376634
rect 564382 376398 582326 376634
rect 582562 376398 582646 376634
rect 582882 376398 586302 376634
rect 586538 376398 586622 376634
rect 586858 376398 592650 376634
rect -8726 376366 592650 376398
rect -8726 372454 592650 372486
rect -8726 372218 -1974 372454
rect -1738 372218 -1654 372454
rect -1418 372218 5826 372454
rect 6062 372218 6146 372454
rect 6382 372218 185826 372454
rect 186062 372218 186146 372454
rect 186382 372218 221826 372454
rect 222062 372218 222146 372454
rect 222382 372218 257826 372454
rect 258062 372218 258146 372454
rect 258382 372218 293826 372454
rect 294062 372218 294146 372454
rect 294382 372218 329826 372454
rect 330062 372218 330146 372454
rect 330382 372218 365826 372454
rect 366062 372218 366146 372454
rect 366382 372218 401826 372454
rect 402062 372218 402146 372454
rect 402382 372218 570350 372454
rect 570586 372218 570670 372454
rect 570906 372218 585342 372454
rect 585578 372218 585662 372454
rect 585898 372218 592650 372454
rect -8726 372134 592650 372218
rect -8726 371898 -1974 372134
rect -1738 371898 -1654 372134
rect -1418 371898 5826 372134
rect 6062 371898 6146 372134
rect 6382 371898 185826 372134
rect 186062 371898 186146 372134
rect 186382 371898 221826 372134
rect 222062 371898 222146 372134
rect 222382 371898 257826 372134
rect 258062 371898 258146 372134
rect 258382 371898 293826 372134
rect 294062 371898 294146 372134
rect 294382 371898 329826 372134
rect 330062 371898 330146 372134
rect 330382 371898 365826 372134
rect 366062 371898 366146 372134
rect 366382 371898 401826 372134
rect 402062 371898 402146 372134
rect 402382 371898 570350 372134
rect 570586 371898 570670 372134
rect 570906 371898 585342 372134
rect 585578 371898 585662 372134
rect 585898 371898 592650 372134
rect -8726 371866 592650 371898
rect -8726 340954 592650 340986
rect -8726 340718 -2934 340954
rect -2698 340718 -2614 340954
rect -2378 340718 13198 340954
rect 13434 340718 13518 340954
rect 13754 340718 167826 340954
rect 168062 340718 168146 340954
rect 168382 340718 203826 340954
rect 204062 340718 204146 340954
rect 204382 340718 239826 340954
rect 240062 340718 240146 340954
rect 240382 340718 275826 340954
rect 276062 340718 276146 340954
rect 276382 340718 311826 340954
rect 312062 340718 312146 340954
rect 312382 340718 347826 340954
rect 348062 340718 348146 340954
rect 348382 340718 383826 340954
rect 384062 340718 384146 340954
rect 384382 340718 419826 340954
rect 420062 340718 420146 340954
rect 420382 340718 563826 340954
rect 564062 340718 564146 340954
rect 564382 340718 582326 340954
rect 582562 340718 582646 340954
rect 582882 340718 586302 340954
rect 586538 340718 586622 340954
rect 586858 340718 592650 340954
rect -8726 340634 592650 340718
rect -8726 340398 -2934 340634
rect -2698 340398 -2614 340634
rect -2378 340398 13198 340634
rect 13434 340398 13518 340634
rect 13754 340398 167826 340634
rect 168062 340398 168146 340634
rect 168382 340398 203826 340634
rect 204062 340398 204146 340634
rect 204382 340398 239826 340634
rect 240062 340398 240146 340634
rect 240382 340398 275826 340634
rect 276062 340398 276146 340634
rect 276382 340398 311826 340634
rect 312062 340398 312146 340634
rect 312382 340398 347826 340634
rect 348062 340398 348146 340634
rect 348382 340398 383826 340634
rect 384062 340398 384146 340634
rect 384382 340398 419826 340634
rect 420062 340398 420146 340634
rect 420382 340398 563826 340634
rect 564062 340398 564146 340634
rect 564382 340398 582326 340634
rect 582562 340398 582646 340634
rect 582882 340398 586302 340634
rect 586538 340398 586622 340634
rect 586858 340398 592650 340634
rect -8726 340366 592650 340398
rect -8726 336454 592650 336486
rect -8726 336218 -1974 336454
rect -1738 336218 -1654 336454
rect -1418 336218 5826 336454
rect 6062 336218 6146 336454
rect 6382 336218 185826 336454
rect 186062 336218 186146 336454
rect 186382 336218 221826 336454
rect 222062 336218 222146 336454
rect 222382 336218 257826 336454
rect 258062 336218 258146 336454
rect 258382 336218 293826 336454
rect 294062 336218 294146 336454
rect 294382 336218 329826 336454
rect 330062 336218 330146 336454
rect 330382 336218 365826 336454
rect 366062 336218 366146 336454
rect 366382 336218 401826 336454
rect 402062 336218 402146 336454
rect 402382 336218 570350 336454
rect 570586 336218 570670 336454
rect 570906 336218 585342 336454
rect 585578 336218 585662 336454
rect 585898 336218 592650 336454
rect -8726 336134 592650 336218
rect -8726 335898 -1974 336134
rect -1738 335898 -1654 336134
rect -1418 335898 5826 336134
rect 6062 335898 6146 336134
rect 6382 335898 185826 336134
rect 186062 335898 186146 336134
rect 186382 335898 221826 336134
rect 222062 335898 222146 336134
rect 222382 335898 257826 336134
rect 258062 335898 258146 336134
rect 258382 335898 293826 336134
rect 294062 335898 294146 336134
rect 294382 335898 329826 336134
rect 330062 335898 330146 336134
rect 330382 335898 365826 336134
rect 366062 335898 366146 336134
rect 366382 335898 401826 336134
rect 402062 335898 402146 336134
rect 402382 335898 570350 336134
rect 570586 335898 570670 336134
rect 570906 335898 585342 336134
rect 585578 335898 585662 336134
rect 585898 335898 592650 336134
rect -8726 335866 592650 335898
rect -8726 304954 592650 304986
rect -8726 304718 -2934 304954
rect -2698 304718 -2614 304954
rect -2378 304718 13198 304954
rect 13434 304718 13518 304954
rect 13754 304718 167826 304954
rect 168062 304718 168146 304954
rect 168382 304718 203826 304954
rect 204062 304718 204146 304954
rect 204382 304718 239826 304954
rect 240062 304718 240146 304954
rect 240382 304718 275826 304954
rect 276062 304718 276146 304954
rect 276382 304718 311826 304954
rect 312062 304718 312146 304954
rect 312382 304718 347826 304954
rect 348062 304718 348146 304954
rect 348382 304718 383826 304954
rect 384062 304718 384146 304954
rect 384382 304718 419826 304954
rect 420062 304718 420146 304954
rect 420382 304718 563826 304954
rect 564062 304718 564146 304954
rect 564382 304718 582326 304954
rect 582562 304718 582646 304954
rect 582882 304718 586302 304954
rect 586538 304718 586622 304954
rect 586858 304718 592650 304954
rect -8726 304634 592650 304718
rect -8726 304398 -2934 304634
rect -2698 304398 -2614 304634
rect -2378 304398 13198 304634
rect 13434 304398 13518 304634
rect 13754 304398 167826 304634
rect 168062 304398 168146 304634
rect 168382 304398 203826 304634
rect 204062 304398 204146 304634
rect 204382 304398 239826 304634
rect 240062 304398 240146 304634
rect 240382 304398 275826 304634
rect 276062 304398 276146 304634
rect 276382 304398 311826 304634
rect 312062 304398 312146 304634
rect 312382 304398 347826 304634
rect 348062 304398 348146 304634
rect 348382 304398 383826 304634
rect 384062 304398 384146 304634
rect 384382 304398 419826 304634
rect 420062 304398 420146 304634
rect 420382 304398 563826 304634
rect 564062 304398 564146 304634
rect 564382 304398 582326 304634
rect 582562 304398 582646 304634
rect 582882 304398 586302 304634
rect 586538 304398 586622 304634
rect 586858 304398 592650 304634
rect -8726 304366 592650 304398
rect -8726 300454 592650 300486
rect -8726 300218 -1974 300454
rect -1738 300218 -1654 300454
rect -1418 300218 5826 300454
rect 6062 300218 6146 300454
rect 6382 300218 185826 300454
rect 186062 300218 186146 300454
rect 186382 300218 221826 300454
rect 222062 300218 222146 300454
rect 222382 300218 257826 300454
rect 258062 300218 258146 300454
rect 258382 300218 293826 300454
rect 294062 300218 294146 300454
rect 294382 300218 329826 300454
rect 330062 300218 330146 300454
rect 330382 300218 365826 300454
rect 366062 300218 366146 300454
rect 366382 300218 401826 300454
rect 402062 300218 402146 300454
rect 402382 300218 570350 300454
rect 570586 300218 570670 300454
rect 570906 300218 585342 300454
rect 585578 300218 585662 300454
rect 585898 300218 592650 300454
rect -8726 300134 592650 300218
rect -8726 299898 -1974 300134
rect -1738 299898 -1654 300134
rect -1418 299898 5826 300134
rect 6062 299898 6146 300134
rect 6382 299898 185826 300134
rect 186062 299898 186146 300134
rect 186382 299898 221826 300134
rect 222062 299898 222146 300134
rect 222382 299898 257826 300134
rect 258062 299898 258146 300134
rect 258382 299898 293826 300134
rect 294062 299898 294146 300134
rect 294382 299898 329826 300134
rect 330062 299898 330146 300134
rect 330382 299898 365826 300134
rect 366062 299898 366146 300134
rect 366382 299898 401826 300134
rect 402062 299898 402146 300134
rect 402382 299898 570350 300134
rect 570586 299898 570670 300134
rect 570906 299898 585342 300134
rect 585578 299898 585662 300134
rect 585898 299898 592650 300134
rect -8726 299866 592650 299898
rect -8726 268954 592650 268986
rect -8726 268718 -2934 268954
rect -2698 268718 -2614 268954
rect -2378 268718 13198 268954
rect 13434 268718 13518 268954
rect 13754 268718 167826 268954
rect 168062 268718 168146 268954
rect 168382 268718 203826 268954
rect 204062 268718 204146 268954
rect 204382 268718 239826 268954
rect 240062 268718 240146 268954
rect 240382 268718 275826 268954
rect 276062 268718 276146 268954
rect 276382 268718 311826 268954
rect 312062 268718 312146 268954
rect 312382 268718 347826 268954
rect 348062 268718 348146 268954
rect 348382 268718 383826 268954
rect 384062 268718 384146 268954
rect 384382 268718 419826 268954
rect 420062 268718 420146 268954
rect 420382 268718 563826 268954
rect 564062 268718 564146 268954
rect 564382 268718 582326 268954
rect 582562 268718 582646 268954
rect 582882 268718 586302 268954
rect 586538 268718 586622 268954
rect 586858 268718 592650 268954
rect -8726 268634 592650 268718
rect -8726 268398 -2934 268634
rect -2698 268398 -2614 268634
rect -2378 268398 13198 268634
rect 13434 268398 13518 268634
rect 13754 268398 167826 268634
rect 168062 268398 168146 268634
rect 168382 268398 203826 268634
rect 204062 268398 204146 268634
rect 204382 268398 239826 268634
rect 240062 268398 240146 268634
rect 240382 268398 275826 268634
rect 276062 268398 276146 268634
rect 276382 268398 311826 268634
rect 312062 268398 312146 268634
rect 312382 268398 347826 268634
rect 348062 268398 348146 268634
rect 348382 268398 383826 268634
rect 384062 268398 384146 268634
rect 384382 268398 419826 268634
rect 420062 268398 420146 268634
rect 420382 268398 563826 268634
rect 564062 268398 564146 268634
rect 564382 268398 582326 268634
rect 582562 268398 582646 268634
rect 582882 268398 586302 268634
rect 586538 268398 586622 268634
rect 586858 268398 592650 268634
rect -8726 268366 592650 268398
rect -8726 264454 592650 264486
rect -8726 264218 -1974 264454
rect -1738 264218 -1654 264454
rect -1418 264218 5826 264454
rect 6062 264218 6146 264454
rect 6382 264218 185826 264454
rect 186062 264218 186146 264454
rect 186382 264218 221826 264454
rect 222062 264218 222146 264454
rect 222382 264218 257826 264454
rect 258062 264218 258146 264454
rect 258382 264218 293826 264454
rect 294062 264218 294146 264454
rect 294382 264218 329826 264454
rect 330062 264218 330146 264454
rect 330382 264218 365826 264454
rect 366062 264218 366146 264454
rect 366382 264218 401826 264454
rect 402062 264218 402146 264454
rect 402382 264218 570350 264454
rect 570586 264218 570670 264454
rect 570906 264218 585342 264454
rect 585578 264218 585662 264454
rect 585898 264218 592650 264454
rect -8726 264134 592650 264218
rect -8726 263898 -1974 264134
rect -1738 263898 -1654 264134
rect -1418 263898 5826 264134
rect 6062 263898 6146 264134
rect 6382 263898 185826 264134
rect 186062 263898 186146 264134
rect 186382 263898 221826 264134
rect 222062 263898 222146 264134
rect 222382 263898 257826 264134
rect 258062 263898 258146 264134
rect 258382 263898 293826 264134
rect 294062 263898 294146 264134
rect 294382 263898 329826 264134
rect 330062 263898 330146 264134
rect 330382 263898 365826 264134
rect 366062 263898 366146 264134
rect 366382 263898 401826 264134
rect 402062 263898 402146 264134
rect 402382 263898 570350 264134
rect 570586 263898 570670 264134
rect 570906 263898 585342 264134
rect 585578 263898 585662 264134
rect 585898 263898 592650 264134
rect -8726 263866 592650 263898
rect -8726 232954 592650 232986
rect -8726 232718 -2934 232954
rect -2698 232718 -2614 232954
rect -2378 232718 23826 232954
rect 24062 232718 24146 232954
rect 24382 232718 59826 232954
rect 60062 232718 60146 232954
rect 60382 232718 95826 232954
rect 96062 232718 96146 232954
rect 96382 232718 131826 232954
rect 132062 232718 132146 232954
rect 132382 232718 167826 232954
rect 168062 232718 168146 232954
rect 168382 232718 203826 232954
rect 204062 232718 204146 232954
rect 204382 232718 239826 232954
rect 240062 232718 240146 232954
rect 240382 232718 275826 232954
rect 276062 232718 276146 232954
rect 276382 232718 311826 232954
rect 312062 232718 312146 232954
rect 312382 232718 347826 232954
rect 348062 232718 348146 232954
rect 348382 232718 383826 232954
rect 384062 232718 384146 232954
rect 384382 232718 419826 232954
rect 420062 232718 420146 232954
rect 420382 232718 455826 232954
rect 456062 232718 456146 232954
rect 456382 232718 491826 232954
rect 492062 232718 492146 232954
rect 492382 232718 527826 232954
rect 528062 232718 528146 232954
rect 528382 232718 563826 232954
rect 564062 232718 564146 232954
rect 564382 232718 582326 232954
rect 582562 232718 582646 232954
rect 582882 232718 586302 232954
rect 586538 232718 586622 232954
rect 586858 232718 592650 232954
rect -8726 232634 592650 232718
rect -8726 232398 -2934 232634
rect -2698 232398 -2614 232634
rect -2378 232398 23826 232634
rect 24062 232398 24146 232634
rect 24382 232398 59826 232634
rect 60062 232398 60146 232634
rect 60382 232398 95826 232634
rect 96062 232398 96146 232634
rect 96382 232398 131826 232634
rect 132062 232398 132146 232634
rect 132382 232398 167826 232634
rect 168062 232398 168146 232634
rect 168382 232398 203826 232634
rect 204062 232398 204146 232634
rect 204382 232398 239826 232634
rect 240062 232398 240146 232634
rect 240382 232398 275826 232634
rect 276062 232398 276146 232634
rect 276382 232398 311826 232634
rect 312062 232398 312146 232634
rect 312382 232398 347826 232634
rect 348062 232398 348146 232634
rect 348382 232398 383826 232634
rect 384062 232398 384146 232634
rect 384382 232398 419826 232634
rect 420062 232398 420146 232634
rect 420382 232398 455826 232634
rect 456062 232398 456146 232634
rect 456382 232398 491826 232634
rect 492062 232398 492146 232634
rect 492382 232398 527826 232634
rect 528062 232398 528146 232634
rect 528382 232398 563826 232634
rect 564062 232398 564146 232634
rect 564382 232398 582326 232634
rect 582562 232398 582646 232634
rect 582882 232398 586302 232634
rect 586538 232398 586622 232634
rect 586858 232398 592650 232634
rect -8726 232366 592650 232398
rect -8726 228454 592650 228486
rect -8726 228218 -1974 228454
rect -1738 228218 -1654 228454
rect -1418 228218 5826 228454
rect 6062 228218 6146 228454
rect 6382 228218 41826 228454
rect 42062 228218 42146 228454
rect 42382 228218 77826 228454
rect 78062 228218 78146 228454
rect 78382 228218 113826 228454
rect 114062 228218 114146 228454
rect 114382 228218 149826 228454
rect 150062 228218 150146 228454
rect 150382 228218 185826 228454
rect 186062 228218 186146 228454
rect 186382 228218 221826 228454
rect 222062 228218 222146 228454
rect 222382 228218 257826 228454
rect 258062 228218 258146 228454
rect 258382 228218 293826 228454
rect 294062 228218 294146 228454
rect 294382 228218 329826 228454
rect 330062 228218 330146 228454
rect 330382 228218 365826 228454
rect 366062 228218 366146 228454
rect 366382 228218 401826 228454
rect 402062 228218 402146 228454
rect 402382 228218 437826 228454
rect 438062 228218 438146 228454
rect 438382 228218 473826 228454
rect 474062 228218 474146 228454
rect 474382 228218 509826 228454
rect 510062 228218 510146 228454
rect 510382 228218 545826 228454
rect 546062 228218 546146 228454
rect 546382 228218 585342 228454
rect 585578 228218 585662 228454
rect 585898 228218 592650 228454
rect -8726 228134 592650 228218
rect -8726 227898 -1974 228134
rect -1738 227898 -1654 228134
rect -1418 227898 5826 228134
rect 6062 227898 6146 228134
rect 6382 227898 41826 228134
rect 42062 227898 42146 228134
rect 42382 227898 77826 228134
rect 78062 227898 78146 228134
rect 78382 227898 113826 228134
rect 114062 227898 114146 228134
rect 114382 227898 149826 228134
rect 150062 227898 150146 228134
rect 150382 227898 185826 228134
rect 186062 227898 186146 228134
rect 186382 227898 221826 228134
rect 222062 227898 222146 228134
rect 222382 227898 257826 228134
rect 258062 227898 258146 228134
rect 258382 227898 293826 228134
rect 294062 227898 294146 228134
rect 294382 227898 329826 228134
rect 330062 227898 330146 228134
rect 330382 227898 365826 228134
rect 366062 227898 366146 228134
rect 366382 227898 401826 228134
rect 402062 227898 402146 228134
rect 402382 227898 437826 228134
rect 438062 227898 438146 228134
rect 438382 227898 473826 228134
rect 474062 227898 474146 228134
rect 474382 227898 509826 228134
rect 510062 227898 510146 228134
rect 510382 227898 545826 228134
rect 546062 227898 546146 228134
rect 546382 227898 585342 228134
rect 585578 227898 585662 228134
rect 585898 227898 592650 228134
rect -8726 227866 592650 227898
rect -8726 196954 592650 196986
rect -8726 196718 -2934 196954
rect -2698 196718 -2614 196954
rect -2378 196718 13198 196954
rect 13434 196718 13518 196954
rect 13754 196718 167826 196954
rect 168062 196718 168146 196954
rect 168382 196718 203826 196954
rect 204062 196718 204146 196954
rect 204382 196718 239826 196954
rect 240062 196718 240146 196954
rect 240382 196718 275826 196954
rect 276062 196718 276146 196954
rect 276382 196718 311826 196954
rect 312062 196718 312146 196954
rect 312382 196718 347826 196954
rect 348062 196718 348146 196954
rect 348382 196718 383826 196954
rect 384062 196718 384146 196954
rect 384382 196718 419826 196954
rect 420062 196718 420146 196954
rect 420382 196718 563826 196954
rect 564062 196718 564146 196954
rect 564382 196718 582326 196954
rect 582562 196718 582646 196954
rect 582882 196718 586302 196954
rect 586538 196718 586622 196954
rect 586858 196718 592650 196954
rect -8726 196634 592650 196718
rect -8726 196398 -2934 196634
rect -2698 196398 -2614 196634
rect -2378 196398 13198 196634
rect 13434 196398 13518 196634
rect 13754 196398 167826 196634
rect 168062 196398 168146 196634
rect 168382 196398 203826 196634
rect 204062 196398 204146 196634
rect 204382 196398 239826 196634
rect 240062 196398 240146 196634
rect 240382 196398 275826 196634
rect 276062 196398 276146 196634
rect 276382 196398 311826 196634
rect 312062 196398 312146 196634
rect 312382 196398 347826 196634
rect 348062 196398 348146 196634
rect 348382 196398 383826 196634
rect 384062 196398 384146 196634
rect 384382 196398 419826 196634
rect 420062 196398 420146 196634
rect 420382 196398 563826 196634
rect 564062 196398 564146 196634
rect 564382 196398 582326 196634
rect 582562 196398 582646 196634
rect 582882 196398 586302 196634
rect 586538 196398 586622 196634
rect 586858 196398 592650 196634
rect -8726 196366 592650 196398
rect -8726 192454 592650 192486
rect -8726 192218 -1974 192454
rect -1738 192218 -1654 192454
rect -1418 192218 5826 192454
rect 6062 192218 6146 192454
rect 6382 192218 185826 192454
rect 186062 192218 186146 192454
rect 186382 192218 221826 192454
rect 222062 192218 222146 192454
rect 222382 192218 257826 192454
rect 258062 192218 258146 192454
rect 258382 192218 293826 192454
rect 294062 192218 294146 192454
rect 294382 192218 329826 192454
rect 330062 192218 330146 192454
rect 330382 192218 365826 192454
rect 366062 192218 366146 192454
rect 366382 192218 401826 192454
rect 402062 192218 402146 192454
rect 402382 192218 570350 192454
rect 570586 192218 570670 192454
rect 570906 192218 585342 192454
rect 585578 192218 585662 192454
rect 585898 192218 592650 192454
rect -8726 192134 592650 192218
rect -8726 191898 -1974 192134
rect -1738 191898 -1654 192134
rect -1418 191898 5826 192134
rect 6062 191898 6146 192134
rect 6382 191898 185826 192134
rect 186062 191898 186146 192134
rect 186382 191898 221826 192134
rect 222062 191898 222146 192134
rect 222382 191898 257826 192134
rect 258062 191898 258146 192134
rect 258382 191898 293826 192134
rect 294062 191898 294146 192134
rect 294382 191898 329826 192134
rect 330062 191898 330146 192134
rect 330382 191898 365826 192134
rect 366062 191898 366146 192134
rect 366382 191898 401826 192134
rect 402062 191898 402146 192134
rect 402382 191898 570350 192134
rect 570586 191898 570670 192134
rect 570906 191898 585342 192134
rect 585578 191898 585662 192134
rect 585898 191898 592650 192134
rect -8726 191866 592650 191898
rect -8726 160954 592650 160986
rect -8726 160718 -2934 160954
rect -2698 160718 -2614 160954
rect -2378 160718 13198 160954
rect 13434 160718 13518 160954
rect 13754 160718 167826 160954
rect 168062 160718 168146 160954
rect 168382 160718 203826 160954
rect 204062 160718 204146 160954
rect 204382 160718 239826 160954
rect 240062 160718 240146 160954
rect 240382 160718 275826 160954
rect 276062 160718 276146 160954
rect 276382 160718 311826 160954
rect 312062 160718 312146 160954
rect 312382 160718 347826 160954
rect 348062 160718 348146 160954
rect 348382 160718 383826 160954
rect 384062 160718 384146 160954
rect 384382 160718 419826 160954
rect 420062 160718 420146 160954
rect 420382 160718 563826 160954
rect 564062 160718 564146 160954
rect 564382 160718 582326 160954
rect 582562 160718 582646 160954
rect 582882 160718 586302 160954
rect 586538 160718 586622 160954
rect 586858 160718 592650 160954
rect -8726 160634 592650 160718
rect -8726 160398 -2934 160634
rect -2698 160398 -2614 160634
rect -2378 160398 13198 160634
rect 13434 160398 13518 160634
rect 13754 160398 167826 160634
rect 168062 160398 168146 160634
rect 168382 160398 203826 160634
rect 204062 160398 204146 160634
rect 204382 160398 239826 160634
rect 240062 160398 240146 160634
rect 240382 160398 275826 160634
rect 276062 160398 276146 160634
rect 276382 160398 311826 160634
rect 312062 160398 312146 160634
rect 312382 160398 347826 160634
rect 348062 160398 348146 160634
rect 348382 160398 383826 160634
rect 384062 160398 384146 160634
rect 384382 160398 419826 160634
rect 420062 160398 420146 160634
rect 420382 160398 563826 160634
rect 564062 160398 564146 160634
rect 564382 160398 582326 160634
rect 582562 160398 582646 160634
rect 582882 160398 586302 160634
rect 586538 160398 586622 160634
rect 586858 160398 592650 160634
rect -8726 160366 592650 160398
rect -8726 156454 592650 156486
rect -8726 156218 -1974 156454
rect -1738 156218 -1654 156454
rect -1418 156218 5826 156454
rect 6062 156218 6146 156454
rect 6382 156218 185826 156454
rect 186062 156218 186146 156454
rect 186382 156218 221826 156454
rect 222062 156218 222146 156454
rect 222382 156218 257826 156454
rect 258062 156218 258146 156454
rect 258382 156218 293826 156454
rect 294062 156218 294146 156454
rect 294382 156218 329826 156454
rect 330062 156218 330146 156454
rect 330382 156218 365826 156454
rect 366062 156218 366146 156454
rect 366382 156218 401826 156454
rect 402062 156218 402146 156454
rect 402382 156218 570350 156454
rect 570586 156218 570670 156454
rect 570906 156218 585342 156454
rect 585578 156218 585662 156454
rect 585898 156218 592650 156454
rect -8726 156134 592650 156218
rect -8726 155898 -1974 156134
rect -1738 155898 -1654 156134
rect -1418 155898 5826 156134
rect 6062 155898 6146 156134
rect 6382 155898 185826 156134
rect 186062 155898 186146 156134
rect 186382 155898 221826 156134
rect 222062 155898 222146 156134
rect 222382 155898 257826 156134
rect 258062 155898 258146 156134
rect 258382 155898 293826 156134
rect 294062 155898 294146 156134
rect 294382 155898 329826 156134
rect 330062 155898 330146 156134
rect 330382 155898 365826 156134
rect 366062 155898 366146 156134
rect 366382 155898 401826 156134
rect 402062 155898 402146 156134
rect 402382 155898 570350 156134
rect 570586 155898 570670 156134
rect 570906 155898 585342 156134
rect 585578 155898 585662 156134
rect 585898 155898 592650 156134
rect -8726 155866 592650 155898
rect -8726 124954 592650 124986
rect -8726 124718 -2934 124954
rect -2698 124718 -2614 124954
rect -2378 124718 23826 124954
rect 24062 124718 24146 124954
rect 24382 124718 59826 124954
rect 60062 124718 60146 124954
rect 60382 124718 95826 124954
rect 96062 124718 96146 124954
rect 96382 124718 131826 124954
rect 132062 124718 132146 124954
rect 132382 124718 167826 124954
rect 168062 124718 168146 124954
rect 168382 124718 203826 124954
rect 204062 124718 204146 124954
rect 204382 124718 239826 124954
rect 240062 124718 240146 124954
rect 240382 124718 275826 124954
rect 276062 124718 276146 124954
rect 276382 124718 311826 124954
rect 312062 124718 312146 124954
rect 312382 124718 347826 124954
rect 348062 124718 348146 124954
rect 348382 124718 383826 124954
rect 384062 124718 384146 124954
rect 384382 124718 419826 124954
rect 420062 124718 420146 124954
rect 420382 124718 455826 124954
rect 456062 124718 456146 124954
rect 456382 124718 491826 124954
rect 492062 124718 492146 124954
rect 492382 124718 527826 124954
rect 528062 124718 528146 124954
rect 528382 124718 563826 124954
rect 564062 124718 564146 124954
rect 564382 124718 582326 124954
rect 582562 124718 582646 124954
rect 582882 124718 586302 124954
rect 586538 124718 586622 124954
rect 586858 124718 592650 124954
rect -8726 124634 592650 124718
rect -8726 124398 -2934 124634
rect -2698 124398 -2614 124634
rect -2378 124398 23826 124634
rect 24062 124398 24146 124634
rect 24382 124398 59826 124634
rect 60062 124398 60146 124634
rect 60382 124398 95826 124634
rect 96062 124398 96146 124634
rect 96382 124398 131826 124634
rect 132062 124398 132146 124634
rect 132382 124398 167826 124634
rect 168062 124398 168146 124634
rect 168382 124398 203826 124634
rect 204062 124398 204146 124634
rect 204382 124398 239826 124634
rect 240062 124398 240146 124634
rect 240382 124398 275826 124634
rect 276062 124398 276146 124634
rect 276382 124398 311826 124634
rect 312062 124398 312146 124634
rect 312382 124398 347826 124634
rect 348062 124398 348146 124634
rect 348382 124398 383826 124634
rect 384062 124398 384146 124634
rect 384382 124398 419826 124634
rect 420062 124398 420146 124634
rect 420382 124398 455826 124634
rect 456062 124398 456146 124634
rect 456382 124398 491826 124634
rect 492062 124398 492146 124634
rect 492382 124398 527826 124634
rect 528062 124398 528146 124634
rect 528382 124398 563826 124634
rect 564062 124398 564146 124634
rect 564382 124398 582326 124634
rect 582562 124398 582646 124634
rect 582882 124398 586302 124634
rect 586538 124398 586622 124634
rect 586858 124398 592650 124634
rect -8726 124366 592650 124398
rect -8726 120454 592650 120486
rect -8726 120218 -1974 120454
rect -1738 120218 -1654 120454
rect -1418 120218 5826 120454
rect 6062 120218 6146 120454
rect 6382 120218 41826 120454
rect 42062 120218 42146 120454
rect 42382 120218 77826 120454
rect 78062 120218 78146 120454
rect 78382 120218 113826 120454
rect 114062 120218 114146 120454
rect 114382 120218 149826 120454
rect 150062 120218 150146 120454
rect 150382 120218 185826 120454
rect 186062 120218 186146 120454
rect 186382 120218 221826 120454
rect 222062 120218 222146 120454
rect 222382 120218 257826 120454
rect 258062 120218 258146 120454
rect 258382 120218 293826 120454
rect 294062 120218 294146 120454
rect 294382 120218 329826 120454
rect 330062 120218 330146 120454
rect 330382 120218 365826 120454
rect 366062 120218 366146 120454
rect 366382 120218 401826 120454
rect 402062 120218 402146 120454
rect 402382 120218 437826 120454
rect 438062 120218 438146 120454
rect 438382 120218 473826 120454
rect 474062 120218 474146 120454
rect 474382 120218 509826 120454
rect 510062 120218 510146 120454
rect 510382 120218 545826 120454
rect 546062 120218 546146 120454
rect 546382 120218 585342 120454
rect 585578 120218 585662 120454
rect 585898 120218 592650 120454
rect -8726 120134 592650 120218
rect -8726 119898 -1974 120134
rect -1738 119898 -1654 120134
rect -1418 119898 5826 120134
rect 6062 119898 6146 120134
rect 6382 119898 41826 120134
rect 42062 119898 42146 120134
rect 42382 119898 77826 120134
rect 78062 119898 78146 120134
rect 78382 119898 113826 120134
rect 114062 119898 114146 120134
rect 114382 119898 149826 120134
rect 150062 119898 150146 120134
rect 150382 119898 185826 120134
rect 186062 119898 186146 120134
rect 186382 119898 221826 120134
rect 222062 119898 222146 120134
rect 222382 119898 257826 120134
rect 258062 119898 258146 120134
rect 258382 119898 293826 120134
rect 294062 119898 294146 120134
rect 294382 119898 329826 120134
rect 330062 119898 330146 120134
rect 330382 119898 365826 120134
rect 366062 119898 366146 120134
rect 366382 119898 401826 120134
rect 402062 119898 402146 120134
rect 402382 119898 437826 120134
rect 438062 119898 438146 120134
rect 438382 119898 473826 120134
rect 474062 119898 474146 120134
rect 474382 119898 509826 120134
rect 510062 119898 510146 120134
rect 510382 119898 545826 120134
rect 546062 119898 546146 120134
rect 546382 119898 585342 120134
rect 585578 119898 585662 120134
rect 585898 119898 592650 120134
rect -8726 119866 592650 119898
rect -8726 88954 592650 88986
rect -8726 88718 -2934 88954
rect -2698 88718 -2614 88954
rect -2378 88718 13198 88954
rect 13434 88718 13518 88954
rect 13754 88718 167826 88954
rect 168062 88718 168146 88954
rect 168382 88718 291590 88954
rect 291826 88718 291910 88954
rect 292146 88718 419826 88954
rect 420062 88718 420146 88954
rect 420382 88718 563826 88954
rect 564062 88718 564146 88954
rect 564382 88718 582326 88954
rect 582562 88718 582646 88954
rect 582882 88718 586302 88954
rect 586538 88718 586622 88954
rect 586858 88718 592650 88954
rect -8726 88634 592650 88718
rect -8726 88398 -2934 88634
rect -2698 88398 -2614 88634
rect -2378 88398 13198 88634
rect 13434 88398 13518 88634
rect 13754 88398 167826 88634
rect 168062 88398 168146 88634
rect 168382 88398 291590 88634
rect 291826 88398 291910 88634
rect 292146 88398 419826 88634
rect 420062 88398 420146 88634
rect 420382 88398 563826 88634
rect 564062 88398 564146 88634
rect 564382 88398 582326 88634
rect 582562 88398 582646 88634
rect 582882 88398 586302 88634
rect 586538 88398 586622 88634
rect 586858 88398 592650 88634
rect -8726 88366 592650 88398
rect -8726 84454 592650 84486
rect -8726 84218 -1974 84454
rect -1738 84218 -1654 84454
rect -1418 84218 5826 84454
rect 6062 84218 6146 84454
rect 6382 84218 173094 84454
rect 173330 84218 173414 84454
rect 173650 84218 293826 84454
rect 294062 84218 294146 84454
rect 294382 84218 401826 84454
rect 402062 84218 402146 84454
rect 402382 84218 570350 84454
rect 570586 84218 570670 84454
rect 570906 84218 585342 84454
rect 585578 84218 585662 84454
rect 585898 84218 592650 84454
rect -8726 84134 592650 84218
rect -8726 83898 -1974 84134
rect -1738 83898 -1654 84134
rect -1418 83898 5826 84134
rect 6062 83898 6146 84134
rect 6382 83898 173094 84134
rect 173330 83898 173414 84134
rect 173650 83898 293826 84134
rect 294062 83898 294146 84134
rect 294382 83898 401826 84134
rect 402062 83898 402146 84134
rect 402382 83898 570350 84134
rect 570586 83898 570670 84134
rect 570906 83898 585342 84134
rect 585578 83898 585662 84134
rect 585898 83898 592650 84134
rect -8726 83866 592650 83898
rect -8726 52954 592650 52986
rect -8726 52718 -2934 52954
rect -2698 52718 -2614 52954
rect -2378 52718 13198 52954
rect 13434 52718 13518 52954
rect 13754 52718 167826 52954
rect 168062 52718 168146 52954
rect 168382 52718 291590 52954
rect 291826 52718 291910 52954
rect 292146 52718 419826 52954
rect 420062 52718 420146 52954
rect 420382 52718 563826 52954
rect 564062 52718 564146 52954
rect 564382 52718 582326 52954
rect 582562 52718 582646 52954
rect 582882 52718 586302 52954
rect 586538 52718 586622 52954
rect 586858 52718 592650 52954
rect -8726 52634 592650 52718
rect -8726 52398 -2934 52634
rect -2698 52398 -2614 52634
rect -2378 52398 13198 52634
rect 13434 52398 13518 52634
rect 13754 52398 167826 52634
rect 168062 52398 168146 52634
rect 168382 52398 291590 52634
rect 291826 52398 291910 52634
rect 292146 52398 419826 52634
rect 420062 52398 420146 52634
rect 420382 52398 563826 52634
rect 564062 52398 564146 52634
rect 564382 52398 582326 52634
rect 582562 52398 582646 52634
rect 582882 52398 586302 52634
rect 586538 52398 586622 52634
rect 586858 52398 592650 52634
rect -8726 52366 592650 52398
rect -8726 48454 592650 48486
rect -8726 48218 -1974 48454
rect -1738 48218 -1654 48454
rect -1418 48218 5826 48454
rect 6062 48218 6146 48454
rect 6382 48218 173094 48454
rect 173330 48218 173414 48454
rect 173650 48218 293826 48454
rect 294062 48218 294146 48454
rect 294382 48218 401826 48454
rect 402062 48218 402146 48454
rect 402382 48218 570350 48454
rect 570586 48218 570670 48454
rect 570906 48218 585342 48454
rect 585578 48218 585662 48454
rect 585898 48218 592650 48454
rect -8726 48134 592650 48218
rect -8726 47898 -1974 48134
rect -1738 47898 -1654 48134
rect -1418 47898 5826 48134
rect 6062 47898 6146 48134
rect 6382 47898 173094 48134
rect 173330 47898 173414 48134
rect 173650 47898 293826 48134
rect 294062 47898 294146 48134
rect 294382 47898 401826 48134
rect 402062 47898 402146 48134
rect 402382 47898 570350 48134
rect 570586 47898 570670 48134
rect 570906 47898 585342 48134
rect 585578 47898 585662 48134
rect 585898 47898 592650 48134
rect -8726 47866 592650 47898
rect -8726 16954 592650 16986
rect -8726 16718 -2934 16954
rect -2698 16718 -2614 16954
rect -2378 16718 23826 16954
rect 24062 16718 24146 16954
rect 24382 16718 59826 16954
rect 60062 16718 60146 16954
rect 60382 16718 95826 16954
rect 96062 16718 96146 16954
rect 96382 16718 131826 16954
rect 132062 16718 132146 16954
rect 132382 16718 167826 16954
rect 168062 16718 168146 16954
rect 168382 16718 203826 16954
rect 204062 16718 204146 16954
rect 204382 16718 239826 16954
rect 240062 16718 240146 16954
rect 240382 16718 275826 16954
rect 276062 16718 276146 16954
rect 276382 16718 311826 16954
rect 312062 16718 312146 16954
rect 312382 16718 347826 16954
rect 348062 16718 348146 16954
rect 348382 16718 383826 16954
rect 384062 16718 384146 16954
rect 384382 16718 419826 16954
rect 420062 16718 420146 16954
rect 420382 16718 455826 16954
rect 456062 16718 456146 16954
rect 456382 16718 491826 16954
rect 492062 16718 492146 16954
rect 492382 16718 527826 16954
rect 528062 16718 528146 16954
rect 528382 16718 563826 16954
rect 564062 16718 564146 16954
rect 564382 16718 582326 16954
rect 582562 16718 582646 16954
rect 582882 16718 586302 16954
rect 586538 16718 586622 16954
rect 586858 16718 592650 16954
rect -8726 16634 592650 16718
rect -8726 16398 -2934 16634
rect -2698 16398 -2614 16634
rect -2378 16398 23826 16634
rect 24062 16398 24146 16634
rect 24382 16398 59826 16634
rect 60062 16398 60146 16634
rect 60382 16398 95826 16634
rect 96062 16398 96146 16634
rect 96382 16398 131826 16634
rect 132062 16398 132146 16634
rect 132382 16398 167826 16634
rect 168062 16398 168146 16634
rect 168382 16398 203826 16634
rect 204062 16398 204146 16634
rect 204382 16398 239826 16634
rect 240062 16398 240146 16634
rect 240382 16398 275826 16634
rect 276062 16398 276146 16634
rect 276382 16398 311826 16634
rect 312062 16398 312146 16634
rect 312382 16398 347826 16634
rect 348062 16398 348146 16634
rect 348382 16398 383826 16634
rect 384062 16398 384146 16634
rect 384382 16398 419826 16634
rect 420062 16398 420146 16634
rect 420382 16398 455826 16634
rect 456062 16398 456146 16634
rect 456382 16398 491826 16634
rect 492062 16398 492146 16634
rect 492382 16398 527826 16634
rect 528062 16398 528146 16634
rect 528382 16398 563826 16634
rect 564062 16398 564146 16634
rect 564382 16398 582326 16634
rect 582562 16398 582646 16634
rect 582882 16398 586302 16634
rect 586538 16398 586622 16634
rect 586858 16398 592650 16634
rect -8726 16366 592650 16398
rect -8726 12454 592650 12486
rect -8726 12218 -1974 12454
rect -1738 12218 -1654 12454
rect -1418 12218 5826 12454
rect 6062 12218 6146 12454
rect 6382 12218 41826 12454
rect 42062 12218 42146 12454
rect 42382 12218 77826 12454
rect 78062 12218 78146 12454
rect 78382 12218 113826 12454
rect 114062 12218 114146 12454
rect 114382 12218 149826 12454
rect 150062 12218 150146 12454
rect 150382 12218 185826 12454
rect 186062 12218 186146 12454
rect 186382 12218 221826 12454
rect 222062 12218 222146 12454
rect 222382 12218 257826 12454
rect 258062 12218 258146 12454
rect 258382 12218 293826 12454
rect 294062 12218 294146 12454
rect 294382 12218 329826 12454
rect 330062 12218 330146 12454
rect 330382 12218 365826 12454
rect 366062 12218 366146 12454
rect 366382 12218 401826 12454
rect 402062 12218 402146 12454
rect 402382 12218 437826 12454
rect 438062 12218 438146 12454
rect 438382 12218 473826 12454
rect 474062 12218 474146 12454
rect 474382 12218 509826 12454
rect 510062 12218 510146 12454
rect 510382 12218 545826 12454
rect 546062 12218 546146 12454
rect 546382 12218 585342 12454
rect 585578 12218 585662 12454
rect 585898 12218 592650 12454
rect -8726 12134 592650 12218
rect -8726 11898 -1974 12134
rect -1738 11898 -1654 12134
rect -1418 11898 5826 12134
rect 6062 11898 6146 12134
rect 6382 11898 41826 12134
rect 42062 11898 42146 12134
rect 42382 11898 77826 12134
rect 78062 11898 78146 12134
rect 78382 11898 113826 12134
rect 114062 11898 114146 12134
rect 114382 11898 149826 12134
rect 150062 11898 150146 12134
rect 150382 11898 185826 12134
rect 186062 11898 186146 12134
rect 186382 11898 221826 12134
rect 222062 11898 222146 12134
rect 222382 11898 257826 12134
rect 258062 11898 258146 12134
rect 258382 11898 293826 12134
rect 294062 11898 294146 12134
rect 294382 11898 329826 12134
rect 330062 11898 330146 12134
rect 330382 11898 365826 12134
rect 366062 11898 366146 12134
rect 366382 11898 401826 12134
rect 402062 11898 402146 12134
rect 402382 11898 437826 12134
rect 438062 11898 438146 12134
rect 438382 11898 473826 12134
rect 474062 11898 474146 12134
rect 474382 11898 509826 12134
rect 510062 11898 510146 12134
rect 510382 11898 545826 12134
rect 546062 11898 546146 12134
rect 546382 11898 585342 12134
rect 585578 11898 585662 12134
rect 585898 11898 592650 12134
rect -8726 11866 592650 11898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 582326 -1306
rect 582562 -1542 582646 -1306
rect 582882 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 582326 -1626
rect 582562 -1862 582646 -1626
rect 582882 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use Marmot  Marmot
timestamp 0
transform 1 0 4000 0 1 4000
box -960 -960 576960 696960
<< labels >>
flabel metal3 s 583520 285276 584960 285516 0 FreeSans 960 0 0 0 analog_io[0]
port 0 nsew signal bidirectional
flabel metal2 s 446098 703520 446210 704960 0 FreeSans 448 90 0 0 analog_io[10]
port 1 nsew signal bidirectional
flabel metal2 s 381146 703520 381258 704960 0 FreeSans 448 90 0 0 analog_io[11]
port 2 nsew signal bidirectional
flabel metal2 s 316286 703520 316398 704960 0 FreeSans 448 90 0 0 analog_io[12]
port 3 nsew signal bidirectional
flabel metal2 s 251426 703520 251538 704960 0 FreeSans 448 90 0 0 analog_io[13]
port 4 nsew signal bidirectional
flabel metal2 s 186474 703520 186586 704960 0 FreeSans 448 90 0 0 analog_io[14]
port 5 nsew signal bidirectional
flabel metal2 s 121614 703520 121726 704960 0 FreeSans 448 90 0 0 analog_io[15]
port 6 nsew signal bidirectional
flabel metal2 s 56754 703520 56866 704960 0 FreeSans 448 90 0 0 analog_io[16]
port 7 nsew signal bidirectional
flabel metal3 s -960 697220 480 697460 0 FreeSans 960 0 0 0 analog_io[17]
port 8 nsew signal bidirectional
flabel metal3 s -960 644996 480 645236 0 FreeSans 960 0 0 0 analog_io[18]
port 9 nsew signal bidirectional
flabel metal3 s -960 592908 480 593148 0 FreeSans 960 0 0 0 analog_io[19]
port 10 nsew signal bidirectional
flabel metal3 s 583520 338452 584960 338692 0 FreeSans 960 0 0 0 analog_io[1]
port 11 nsew signal bidirectional
flabel metal3 s -960 540684 480 540924 0 FreeSans 960 0 0 0 analog_io[20]
port 12 nsew signal bidirectional
flabel metal3 s -960 488596 480 488836 0 FreeSans 960 0 0 0 analog_io[21]
port 13 nsew signal bidirectional
flabel metal3 s -960 436508 480 436748 0 FreeSans 960 0 0 0 analog_io[22]
port 14 nsew signal bidirectional
flabel metal3 s -960 384284 480 384524 0 FreeSans 960 0 0 0 analog_io[23]
port 15 nsew signal bidirectional
flabel metal3 s -960 332196 480 332436 0 FreeSans 960 0 0 0 analog_io[24]
port 16 nsew signal bidirectional
flabel metal3 s -960 279972 480 280212 0 FreeSans 960 0 0 0 analog_io[25]
port 17 nsew signal bidirectional
flabel metal3 s -960 227884 480 228124 0 FreeSans 960 0 0 0 analog_io[26]
port 18 nsew signal bidirectional
flabel metal3 s -960 175796 480 176036 0 FreeSans 960 0 0 0 analog_io[27]
port 19 nsew signal bidirectional
flabel metal3 s -960 123572 480 123812 0 FreeSans 960 0 0 0 analog_io[28]
port 20 nsew signal bidirectional
flabel metal3 s 583520 391628 584960 391868 0 FreeSans 960 0 0 0 analog_io[2]
port 21 nsew signal bidirectional
flabel metal3 s 583520 444668 584960 444908 0 FreeSans 960 0 0 0 analog_io[3]
port 22 nsew signal bidirectional
flabel metal3 s 583520 497844 584960 498084 0 FreeSans 960 0 0 0 analog_io[4]
port 23 nsew signal bidirectional
flabel metal3 s 583520 551020 584960 551260 0 FreeSans 960 0 0 0 analog_io[5]
port 24 nsew signal bidirectional
flabel metal3 s 583520 604060 584960 604300 0 FreeSans 960 0 0 0 analog_io[6]
port 25 nsew signal bidirectional
flabel metal3 s 583520 657236 584960 657476 0 FreeSans 960 0 0 0 analog_io[7]
port 26 nsew signal bidirectional
flabel metal2 s 575818 703520 575930 704960 0 FreeSans 448 90 0 0 analog_io[8]
port 27 nsew signal bidirectional
flabel metal2 s 510958 703520 511070 704960 0 FreeSans 448 90 0 0 analog_io[9]
port 28 nsew signal bidirectional
flabel metal3 s 583520 6476 584960 6716 0 FreeSans 960 0 0 0 io_in[0]
port 29 nsew signal input
flabel metal3 s 583520 457996 584960 458236 0 FreeSans 960 0 0 0 io_in[10]
port 30 nsew signal input
flabel metal3 s 583520 511172 584960 511412 0 FreeSans 960 0 0 0 io_in[11]
port 31 nsew signal input
flabel metal3 s 583520 564212 584960 564452 0 FreeSans 960 0 0 0 io_in[12]
port 32 nsew signal input
flabel metal3 s 583520 617388 584960 617628 0 FreeSans 960 0 0 0 io_in[13]
port 33 nsew signal input
flabel metal3 s 583520 670564 584960 670804 0 FreeSans 960 0 0 0 io_in[14]
port 34 nsew signal input
flabel metal2 s 559626 703520 559738 704960 0 FreeSans 448 90 0 0 io_in[15]
port 35 nsew signal input
flabel metal2 s 494766 703520 494878 704960 0 FreeSans 448 90 0 0 io_in[16]
port 36 nsew signal input
flabel metal2 s 429814 703520 429926 704960 0 FreeSans 448 90 0 0 io_in[17]
port 37 nsew signal input
flabel metal2 s 364954 703520 365066 704960 0 FreeSans 448 90 0 0 io_in[18]
port 38 nsew signal input
flabel metal2 s 300094 703520 300206 704960 0 FreeSans 448 90 0 0 io_in[19]
port 39 nsew signal input
flabel metal3 s 583520 46188 584960 46428 0 FreeSans 960 0 0 0 io_in[1]
port 40 nsew signal input
flabel metal2 s 235142 703520 235254 704960 0 FreeSans 448 90 0 0 io_in[20]
port 41 nsew signal input
flabel metal2 s 170282 703520 170394 704960 0 FreeSans 448 90 0 0 io_in[21]
port 42 nsew signal input
flabel metal2 s 105422 703520 105534 704960 0 FreeSans 448 90 0 0 io_in[22]
port 43 nsew signal input
flabel metal2 s 40470 703520 40582 704960 0 FreeSans 448 90 0 0 io_in[23]
port 44 nsew signal input
flabel metal3 s -960 684164 480 684404 0 FreeSans 960 0 0 0 io_in[24]
port 45 nsew signal input
flabel metal3 s -960 631940 480 632180 0 FreeSans 960 0 0 0 io_in[25]
port 46 nsew signal input
flabel metal3 s -960 579852 480 580092 0 FreeSans 960 0 0 0 io_in[26]
port 47 nsew signal input
flabel metal3 s -960 527764 480 528004 0 FreeSans 960 0 0 0 io_in[27]
port 48 nsew signal input
flabel metal3 s -960 475540 480 475780 0 FreeSans 960 0 0 0 io_in[28]
port 49 nsew signal input
flabel metal3 s -960 423452 480 423692 0 FreeSans 960 0 0 0 io_in[29]
port 50 nsew signal input
flabel metal3 s 583520 86036 584960 86276 0 FreeSans 960 0 0 0 io_in[2]
port 51 nsew signal input
flabel metal3 s -960 371228 480 371468 0 FreeSans 960 0 0 0 io_in[30]
port 52 nsew signal input
flabel metal3 s -960 319140 480 319380 0 FreeSans 960 0 0 0 io_in[31]
port 53 nsew signal input
flabel metal3 s -960 267052 480 267292 0 FreeSans 960 0 0 0 io_in[32]
port 54 nsew signal input
flabel metal3 s -960 214828 480 215068 0 FreeSans 960 0 0 0 io_in[33]
port 55 nsew signal input
flabel metal3 s -960 162740 480 162980 0 FreeSans 960 0 0 0 io_in[34]
port 56 nsew signal input
flabel metal3 s -960 110516 480 110756 0 FreeSans 960 0 0 0 io_in[35]
port 57 nsew signal input
flabel metal3 s -960 71484 480 71724 0 FreeSans 960 0 0 0 io_in[36]
port 58 nsew signal input
flabel metal3 s -960 32316 480 32556 0 FreeSans 960 0 0 0 io_in[37]
port 59 nsew signal input
flabel metal3 s 583520 125884 584960 126124 0 FreeSans 960 0 0 0 io_in[3]
port 60 nsew signal input
flabel metal3 s 583520 165732 584960 165972 0 FreeSans 960 0 0 0 io_in[4]
port 61 nsew signal input
flabel metal3 s 583520 205580 584960 205820 0 FreeSans 960 0 0 0 io_in[5]
port 62 nsew signal input
flabel metal3 s 583520 245428 584960 245668 0 FreeSans 960 0 0 0 io_in[6]
port 63 nsew signal input
flabel metal3 s 583520 298604 584960 298844 0 FreeSans 960 0 0 0 io_in[7]
port 64 nsew signal input
flabel metal3 s 583520 351780 584960 352020 0 FreeSans 960 0 0 0 io_in[8]
port 65 nsew signal input
flabel metal3 s 583520 404820 584960 405060 0 FreeSans 960 0 0 0 io_in[9]
port 66 nsew signal input
flabel metal3 s 583520 32996 584960 33236 0 FreeSans 960 0 0 0 io_oeb[0]
port 67 nsew signal tristate
flabel metal3 s 583520 484516 584960 484756 0 FreeSans 960 0 0 0 io_oeb[10]
port 68 nsew signal tristate
flabel metal3 s 583520 537692 584960 537932 0 FreeSans 960 0 0 0 io_oeb[11]
port 69 nsew signal tristate
flabel metal3 s 583520 590868 584960 591108 0 FreeSans 960 0 0 0 io_oeb[12]
port 70 nsew signal tristate
flabel metal3 s 583520 643908 584960 644148 0 FreeSans 960 0 0 0 io_oeb[13]
port 71 nsew signal tristate
flabel metal3 s 583520 697084 584960 697324 0 FreeSans 960 0 0 0 io_oeb[14]
port 72 nsew signal tristate
flabel metal2 s 527150 703520 527262 704960 0 FreeSans 448 90 0 0 io_oeb[15]
port 73 nsew signal tristate
flabel metal2 s 462290 703520 462402 704960 0 FreeSans 448 90 0 0 io_oeb[16]
port 74 nsew signal tristate
flabel metal2 s 397430 703520 397542 704960 0 FreeSans 448 90 0 0 io_oeb[17]
port 75 nsew signal tristate
flabel metal2 s 332478 703520 332590 704960 0 FreeSans 448 90 0 0 io_oeb[18]
port 76 nsew signal tristate
flabel metal2 s 267618 703520 267730 704960 0 FreeSans 448 90 0 0 io_oeb[19]
port 77 nsew signal tristate
flabel metal3 s 583520 72844 584960 73084 0 FreeSans 960 0 0 0 io_oeb[1]
port 78 nsew signal tristate
flabel metal2 s 202758 703520 202870 704960 0 FreeSans 448 90 0 0 io_oeb[20]
port 79 nsew signal tristate
flabel metal2 s 137806 703520 137918 704960 0 FreeSans 448 90 0 0 io_oeb[21]
port 80 nsew signal tristate
flabel metal2 s 72946 703520 73058 704960 0 FreeSans 448 90 0 0 io_oeb[22]
port 81 nsew signal tristate
flabel metal2 s 8086 703520 8198 704960 0 FreeSans 448 90 0 0 io_oeb[23]
port 82 nsew signal tristate
flabel metal3 s -960 658052 480 658292 0 FreeSans 960 0 0 0 io_oeb[24]
port 83 nsew signal tristate
flabel metal3 s -960 605964 480 606204 0 FreeSans 960 0 0 0 io_oeb[25]
port 84 nsew signal tristate
flabel metal3 s -960 553740 480 553980 0 FreeSans 960 0 0 0 io_oeb[26]
port 85 nsew signal tristate
flabel metal3 s -960 501652 480 501892 0 FreeSans 960 0 0 0 io_oeb[27]
port 86 nsew signal tristate
flabel metal3 s -960 449428 480 449668 0 FreeSans 960 0 0 0 io_oeb[28]
port 87 nsew signal tristate
flabel metal3 s -960 397340 480 397580 0 FreeSans 960 0 0 0 io_oeb[29]
port 88 nsew signal tristate
flabel metal3 s 583520 112692 584960 112932 0 FreeSans 960 0 0 0 io_oeb[2]
port 89 nsew signal tristate
flabel metal3 s -960 345252 480 345492 0 FreeSans 960 0 0 0 io_oeb[30]
port 90 nsew signal tristate
flabel metal3 s -960 293028 480 293268 0 FreeSans 960 0 0 0 io_oeb[31]
port 91 nsew signal tristate
flabel metal3 s -960 240940 480 241180 0 FreeSans 960 0 0 0 io_oeb[32]
port 92 nsew signal tristate
flabel metal3 s -960 188716 480 188956 0 FreeSans 960 0 0 0 io_oeb[33]
port 93 nsew signal tristate
flabel metal3 s -960 136628 480 136868 0 FreeSans 960 0 0 0 io_oeb[34]
port 94 nsew signal tristate
flabel metal3 s -960 84540 480 84780 0 FreeSans 960 0 0 0 io_oeb[35]
port 95 nsew signal tristate
flabel metal3 s -960 45372 480 45612 0 FreeSans 960 0 0 0 io_oeb[36]
port 96 nsew signal tristate
flabel metal3 s -960 6340 480 6580 0 FreeSans 960 0 0 0 io_oeb[37]
port 97 nsew signal tristate
flabel metal3 s 583520 152540 584960 152780 0 FreeSans 960 0 0 0 io_oeb[3]
port 98 nsew signal tristate
flabel metal3 s 583520 192388 584960 192628 0 FreeSans 960 0 0 0 io_oeb[4]
port 99 nsew signal tristate
flabel metal3 s 583520 232236 584960 232476 0 FreeSans 960 0 0 0 io_oeb[5]
port 100 nsew signal tristate
flabel metal3 s 583520 272084 584960 272324 0 FreeSans 960 0 0 0 io_oeb[6]
port 101 nsew signal tristate
flabel metal3 s 583520 325124 584960 325364 0 FreeSans 960 0 0 0 io_oeb[7]
port 102 nsew signal tristate
flabel metal3 s 583520 378300 584960 378540 0 FreeSans 960 0 0 0 io_oeb[8]
port 103 nsew signal tristate
flabel metal3 s 583520 431476 584960 431716 0 FreeSans 960 0 0 0 io_oeb[9]
port 104 nsew signal tristate
flabel metal3 s 583520 19668 584960 19908 0 FreeSans 960 0 0 0 io_out[0]
port 105 nsew signal tristate
flabel metal3 s 583520 471324 584960 471564 0 FreeSans 960 0 0 0 io_out[10]
port 106 nsew signal tristate
flabel metal3 s 583520 524364 584960 524604 0 FreeSans 960 0 0 0 io_out[11]
port 107 nsew signal tristate
flabel metal3 s 583520 577540 584960 577780 0 FreeSans 960 0 0 0 io_out[12]
port 108 nsew signal tristate
flabel metal3 s 583520 630716 584960 630956 0 FreeSans 960 0 0 0 io_out[13]
port 109 nsew signal tristate
flabel metal3 s 583520 683756 584960 683996 0 FreeSans 960 0 0 0 io_out[14]
port 110 nsew signal tristate
flabel metal2 s 543434 703520 543546 704960 0 FreeSans 448 90 0 0 io_out[15]
port 111 nsew signal tristate
flabel metal2 s 478482 703520 478594 704960 0 FreeSans 448 90 0 0 io_out[16]
port 112 nsew signal tristate
flabel metal2 s 413622 703520 413734 704960 0 FreeSans 448 90 0 0 io_out[17]
port 113 nsew signal tristate
flabel metal2 s 348762 703520 348874 704960 0 FreeSans 448 90 0 0 io_out[18]
port 114 nsew signal tristate
flabel metal2 s 283810 703520 283922 704960 0 FreeSans 448 90 0 0 io_out[19]
port 115 nsew signal tristate
flabel metal3 s 583520 59516 584960 59756 0 FreeSans 960 0 0 0 io_out[1]
port 116 nsew signal tristate
flabel metal2 s 218950 703520 219062 704960 0 FreeSans 448 90 0 0 io_out[20]
port 117 nsew signal tristate
flabel metal2 s 154090 703520 154202 704960 0 FreeSans 448 90 0 0 io_out[21]
port 118 nsew signal tristate
flabel metal2 s 89138 703520 89250 704960 0 FreeSans 448 90 0 0 io_out[22]
port 119 nsew signal tristate
flabel metal2 s 24278 703520 24390 704960 0 FreeSans 448 90 0 0 io_out[23]
port 120 nsew signal tristate
flabel metal3 s -960 671108 480 671348 0 FreeSans 960 0 0 0 io_out[24]
port 121 nsew signal tristate
flabel metal3 s -960 619020 480 619260 0 FreeSans 960 0 0 0 io_out[25]
port 122 nsew signal tristate
flabel metal3 s -960 566796 480 567036 0 FreeSans 960 0 0 0 io_out[26]
port 123 nsew signal tristate
flabel metal3 s -960 514708 480 514948 0 FreeSans 960 0 0 0 io_out[27]
port 124 nsew signal tristate
flabel metal3 s -960 462484 480 462724 0 FreeSans 960 0 0 0 io_out[28]
port 125 nsew signal tristate
flabel metal3 s -960 410396 480 410636 0 FreeSans 960 0 0 0 io_out[29]
port 126 nsew signal tristate
flabel metal3 s 583520 99364 584960 99604 0 FreeSans 960 0 0 0 io_out[2]
port 127 nsew signal tristate
flabel metal3 s -960 358308 480 358548 0 FreeSans 960 0 0 0 io_out[30]
port 128 nsew signal tristate
flabel metal3 s -960 306084 480 306324 0 FreeSans 960 0 0 0 io_out[31]
port 129 nsew signal tristate
flabel metal3 s -960 253996 480 254236 0 FreeSans 960 0 0 0 io_out[32]
port 130 nsew signal tristate
flabel metal3 s -960 201772 480 202012 0 FreeSans 960 0 0 0 io_out[33]
port 131 nsew signal tristate
flabel metal3 s -960 149684 480 149924 0 FreeSans 960 0 0 0 io_out[34]
port 132 nsew signal tristate
flabel metal3 s -960 97460 480 97700 0 FreeSans 960 0 0 0 io_out[35]
port 133 nsew signal tristate
flabel metal3 s -960 58428 480 58668 0 FreeSans 960 0 0 0 io_out[36]
port 134 nsew signal tristate
flabel metal3 s -960 19260 480 19500 0 FreeSans 960 0 0 0 io_out[37]
port 135 nsew signal tristate
flabel metal3 s 583520 139212 584960 139452 0 FreeSans 960 0 0 0 io_out[3]
port 136 nsew signal tristate
flabel metal3 s 583520 179060 584960 179300 0 FreeSans 960 0 0 0 io_out[4]
port 137 nsew signal tristate
flabel metal3 s 583520 218908 584960 219148 0 FreeSans 960 0 0 0 io_out[5]
port 138 nsew signal tristate
flabel metal3 s 583520 258756 584960 258996 0 FreeSans 960 0 0 0 io_out[6]
port 139 nsew signal tristate
flabel metal3 s 583520 311932 584960 312172 0 FreeSans 960 0 0 0 io_out[7]
port 140 nsew signal tristate
flabel metal3 s 583520 364972 584960 365212 0 FreeSans 960 0 0 0 io_out[8]
port 141 nsew signal tristate
flabel metal3 s 583520 418148 584960 418388 0 FreeSans 960 0 0 0 io_out[9]
port 142 nsew signal tristate
flabel metal2 s 125846 -960 125958 480 0 FreeSans 448 90 0 0 la_data_in[0]
port 143 nsew signal input
flabel metal2 s 480506 -960 480618 480 0 FreeSans 448 90 0 0 la_data_in[100]
port 144 nsew signal input
flabel metal2 s 484002 -960 484114 480 0 FreeSans 448 90 0 0 la_data_in[101]
port 145 nsew signal input
flabel metal2 s 487590 -960 487702 480 0 FreeSans 448 90 0 0 la_data_in[102]
port 146 nsew signal input
flabel metal2 s 491086 -960 491198 480 0 FreeSans 448 90 0 0 la_data_in[103]
port 147 nsew signal input
flabel metal2 s 494674 -960 494786 480 0 FreeSans 448 90 0 0 la_data_in[104]
port 148 nsew signal input
flabel metal2 s 498170 -960 498282 480 0 FreeSans 448 90 0 0 la_data_in[105]
port 149 nsew signal input
flabel metal2 s 501758 -960 501870 480 0 FreeSans 448 90 0 0 la_data_in[106]
port 150 nsew signal input
flabel metal2 s 505346 -960 505458 480 0 FreeSans 448 90 0 0 la_data_in[107]
port 151 nsew signal input
flabel metal2 s 508842 -960 508954 480 0 FreeSans 448 90 0 0 la_data_in[108]
port 152 nsew signal input
flabel metal2 s 512430 -960 512542 480 0 FreeSans 448 90 0 0 la_data_in[109]
port 153 nsew signal input
flabel metal2 s 161266 -960 161378 480 0 FreeSans 448 90 0 0 la_data_in[10]
port 154 nsew signal input
flabel metal2 s 515926 -960 516038 480 0 FreeSans 448 90 0 0 la_data_in[110]
port 155 nsew signal input
flabel metal2 s 519514 -960 519626 480 0 FreeSans 448 90 0 0 la_data_in[111]
port 156 nsew signal input
flabel metal2 s 523010 -960 523122 480 0 FreeSans 448 90 0 0 la_data_in[112]
port 157 nsew signal input
flabel metal2 s 526598 -960 526710 480 0 FreeSans 448 90 0 0 la_data_in[113]
port 158 nsew signal input
flabel metal2 s 530094 -960 530206 480 0 FreeSans 448 90 0 0 la_data_in[114]
port 159 nsew signal input
flabel metal2 s 533682 -960 533794 480 0 FreeSans 448 90 0 0 la_data_in[115]
port 160 nsew signal input
flabel metal2 s 537178 -960 537290 480 0 FreeSans 448 90 0 0 la_data_in[116]
port 161 nsew signal input
flabel metal2 s 540766 -960 540878 480 0 FreeSans 448 90 0 0 la_data_in[117]
port 162 nsew signal input
flabel metal2 s 544354 -960 544466 480 0 FreeSans 448 90 0 0 la_data_in[118]
port 163 nsew signal input
flabel metal2 s 547850 -960 547962 480 0 FreeSans 448 90 0 0 la_data_in[119]
port 164 nsew signal input
flabel metal2 s 164854 -960 164966 480 0 FreeSans 448 90 0 0 la_data_in[11]
port 165 nsew signal input
flabel metal2 s 551438 -960 551550 480 0 FreeSans 448 90 0 0 la_data_in[120]
port 166 nsew signal input
flabel metal2 s 554934 -960 555046 480 0 FreeSans 448 90 0 0 la_data_in[121]
port 167 nsew signal input
flabel metal2 s 558522 -960 558634 480 0 FreeSans 448 90 0 0 la_data_in[122]
port 168 nsew signal input
flabel metal2 s 562018 -960 562130 480 0 FreeSans 448 90 0 0 la_data_in[123]
port 169 nsew signal input
flabel metal2 s 565606 -960 565718 480 0 FreeSans 448 90 0 0 la_data_in[124]
port 170 nsew signal input
flabel metal2 s 569102 -960 569214 480 0 FreeSans 448 90 0 0 la_data_in[125]
port 171 nsew signal input
flabel metal2 s 572690 -960 572802 480 0 FreeSans 448 90 0 0 la_data_in[126]
port 172 nsew signal input
flabel metal2 s 576278 -960 576390 480 0 FreeSans 448 90 0 0 la_data_in[127]
port 173 nsew signal input
flabel metal2 s 168350 -960 168462 480 0 FreeSans 448 90 0 0 la_data_in[12]
port 174 nsew signal input
flabel metal2 s 171938 -960 172050 480 0 FreeSans 448 90 0 0 la_data_in[13]
port 175 nsew signal input
flabel metal2 s 175434 -960 175546 480 0 FreeSans 448 90 0 0 la_data_in[14]
port 176 nsew signal input
flabel metal2 s 179022 -960 179134 480 0 FreeSans 448 90 0 0 la_data_in[15]
port 177 nsew signal input
flabel metal2 s 182518 -960 182630 480 0 FreeSans 448 90 0 0 la_data_in[16]
port 178 nsew signal input
flabel metal2 s 186106 -960 186218 480 0 FreeSans 448 90 0 0 la_data_in[17]
port 179 nsew signal input
flabel metal2 s 189694 -960 189806 480 0 FreeSans 448 90 0 0 la_data_in[18]
port 180 nsew signal input
flabel metal2 s 193190 -960 193302 480 0 FreeSans 448 90 0 0 la_data_in[19]
port 181 nsew signal input
flabel metal2 s 129342 -960 129454 480 0 FreeSans 448 90 0 0 la_data_in[1]
port 182 nsew signal input
flabel metal2 s 196778 -960 196890 480 0 FreeSans 448 90 0 0 la_data_in[20]
port 183 nsew signal input
flabel metal2 s 200274 -960 200386 480 0 FreeSans 448 90 0 0 la_data_in[21]
port 184 nsew signal input
flabel metal2 s 203862 -960 203974 480 0 FreeSans 448 90 0 0 la_data_in[22]
port 185 nsew signal input
flabel metal2 s 207358 -960 207470 480 0 FreeSans 448 90 0 0 la_data_in[23]
port 186 nsew signal input
flabel metal2 s 210946 -960 211058 480 0 FreeSans 448 90 0 0 la_data_in[24]
port 187 nsew signal input
flabel metal2 s 214442 -960 214554 480 0 FreeSans 448 90 0 0 la_data_in[25]
port 188 nsew signal input
flabel metal2 s 218030 -960 218142 480 0 FreeSans 448 90 0 0 la_data_in[26]
port 189 nsew signal input
flabel metal2 s 221526 -960 221638 480 0 FreeSans 448 90 0 0 la_data_in[27]
port 190 nsew signal input
flabel metal2 s 225114 -960 225226 480 0 FreeSans 448 90 0 0 la_data_in[28]
port 191 nsew signal input
flabel metal2 s 228702 -960 228814 480 0 FreeSans 448 90 0 0 la_data_in[29]
port 192 nsew signal input
flabel metal2 s 132930 -960 133042 480 0 FreeSans 448 90 0 0 la_data_in[2]
port 193 nsew signal input
flabel metal2 s 232198 -960 232310 480 0 FreeSans 448 90 0 0 la_data_in[30]
port 194 nsew signal input
flabel metal2 s 235786 -960 235898 480 0 FreeSans 448 90 0 0 la_data_in[31]
port 195 nsew signal input
flabel metal2 s 239282 -960 239394 480 0 FreeSans 448 90 0 0 la_data_in[32]
port 196 nsew signal input
flabel metal2 s 242870 -960 242982 480 0 FreeSans 448 90 0 0 la_data_in[33]
port 197 nsew signal input
flabel metal2 s 246366 -960 246478 480 0 FreeSans 448 90 0 0 la_data_in[34]
port 198 nsew signal input
flabel metal2 s 249954 -960 250066 480 0 FreeSans 448 90 0 0 la_data_in[35]
port 199 nsew signal input
flabel metal2 s 253450 -960 253562 480 0 FreeSans 448 90 0 0 la_data_in[36]
port 200 nsew signal input
flabel metal2 s 257038 -960 257150 480 0 FreeSans 448 90 0 0 la_data_in[37]
port 201 nsew signal input
flabel metal2 s 260626 -960 260738 480 0 FreeSans 448 90 0 0 la_data_in[38]
port 202 nsew signal input
flabel metal2 s 264122 -960 264234 480 0 FreeSans 448 90 0 0 la_data_in[39]
port 203 nsew signal input
flabel metal2 s 136426 -960 136538 480 0 FreeSans 448 90 0 0 la_data_in[3]
port 204 nsew signal input
flabel metal2 s 267710 -960 267822 480 0 FreeSans 448 90 0 0 la_data_in[40]
port 205 nsew signal input
flabel metal2 s 271206 -960 271318 480 0 FreeSans 448 90 0 0 la_data_in[41]
port 206 nsew signal input
flabel metal2 s 274794 -960 274906 480 0 FreeSans 448 90 0 0 la_data_in[42]
port 207 nsew signal input
flabel metal2 s 278290 -960 278402 480 0 FreeSans 448 90 0 0 la_data_in[43]
port 208 nsew signal input
flabel metal2 s 281878 -960 281990 480 0 FreeSans 448 90 0 0 la_data_in[44]
port 209 nsew signal input
flabel metal2 s 285374 -960 285486 480 0 FreeSans 448 90 0 0 la_data_in[45]
port 210 nsew signal input
flabel metal2 s 288962 -960 289074 480 0 FreeSans 448 90 0 0 la_data_in[46]
port 211 nsew signal input
flabel metal2 s 292550 -960 292662 480 0 FreeSans 448 90 0 0 la_data_in[47]
port 212 nsew signal input
flabel metal2 s 296046 -960 296158 480 0 FreeSans 448 90 0 0 la_data_in[48]
port 213 nsew signal input
flabel metal2 s 299634 -960 299746 480 0 FreeSans 448 90 0 0 la_data_in[49]
port 214 nsew signal input
flabel metal2 s 140014 -960 140126 480 0 FreeSans 448 90 0 0 la_data_in[4]
port 215 nsew signal input
flabel metal2 s 303130 -960 303242 480 0 FreeSans 448 90 0 0 la_data_in[50]
port 216 nsew signal input
flabel metal2 s 306718 -960 306830 480 0 FreeSans 448 90 0 0 la_data_in[51]
port 217 nsew signal input
flabel metal2 s 310214 -960 310326 480 0 FreeSans 448 90 0 0 la_data_in[52]
port 218 nsew signal input
flabel metal2 s 313802 -960 313914 480 0 FreeSans 448 90 0 0 la_data_in[53]
port 219 nsew signal input
flabel metal2 s 317298 -960 317410 480 0 FreeSans 448 90 0 0 la_data_in[54]
port 220 nsew signal input
flabel metal2 s 320886 -960 320998 480 0 FreeSans 448 90 0 0 la_data_in[55]
port 221 nsew signal input
flabel metal2 s 324382 -960 324494 480 0 FreeSans 448 90 0 0 la_data_in[56]
port 222 nsew signal input
flabel metal2 s 327970 -960 328082 480 0 FreeSans 448 90 0 0 la_data_in[57]
port 223 nsew signal input
flabel metal2 s 331558 -960 331670 480 0 FreeSans 448 90 0 0 la_data_in[58]
port 224 nsew signal input
flabel metal2 s 335054 -960 335166 480 0 FreeSans 448 90 0 0 la_data_in[59]
port 225 nsew signal input
flabel metal2 s 143510 -960 143622 480 0 FreeSans 448 90 0 0 la_data_in[5]
port 226 nsew signal input
flabel metal2 s 338642 -960 338754 480 0 FreeSans 448 90 0 0 la_data_in[60]
port 227 nsew signal input
flabel metal2 s 342138 -960 342250 480 0 FreeSans 448 90 0 0 la_data_in[61]
port 228 nsew signal input
flabel metal2 s 345726 -960 345838 480 0 FreeSans 448 90 0 0 la_data_in[62]
port 229 nsew signal input
flabel metal2 s 349222 -960 349334 480 0 FreeSans 448 90 0 0 la_data_in[63]
port 230 nsew signal input
flabel metal2 s 352810 -960 352922 480 0 FreeSans 448 90 0 0 la_data_in[64]
port 231 nsew signal input
flabel metal2 s 356306 -960 356418 480 0 FreeSans 448 90 0 0 la_data_in[65]
port 232 nsew signal input
flabel metal2 s 359894 -960 360006 480 0 FreeSans 448 90 0 0 la_data_in[66]
port 233 nsew signal input
flabel metal2 s 363482 -960 363594 480 0 FreeSans 448 90 0 0 la_data_in[67]
port 234 nsew signal input
flabel metal2 s 366978 -960 367090 480 0 FreeSans 448 90 0 0 la_data_in[68]
port 235 nsew signal input
flabel metal2 s 370566 -960 370678 480 0 FreeSans 448 90 0 0 la_data_in[69]
port 236 nsew signal input
flabel metal2 s 147098 -960 147210 480 0 FreeSans 448 90 0 0 la_data_in[6]
port 237 nsew signal input
flabel metal2 s 374062 -960 374174 480 0 FreeSans 448 90 0 0 la_data_in[70]
port 238 nsew signal input
flabel metal2 s 377650 -960 377762 480 0 FreeSans 448 90 0 0 la_data_in[71]
port 239 nsew signal input
flabel metal2 s 381146 -960 381258 480 0 FreeSans 448 90 0 0 la_data_in[72]
port 240 nsew signal input
flabel metal2 s 384734 -960 384846 480 0 FreeSans 448 90 0 0 la_data_in[73]
port 241 nsew signal input
flabel metal2 s 388230 -960 388342 480 0 FreeSans 448 90 0 0 la_data_in[74]
port 242 nsew signal input
flabel metal2 s 391818 -960 391930 480 0 FreeSans 448 90 0 0 la_data_in[75]
port 243 nsew signal input
flabel metal2 s 395314 -960 395426 480 0 FreeSans 448 90 0 0 la_data_in[76]
port 244 nsew signal input
flabel metal2 s 398902 -960 399014 480 0 FreeSans 448 90 0 0 la_data_in[77]
port 245 nsew signal input
flabel metal2 s 402490 -960 402602 480 0 FreeSans 448 90 0 0 la_data_in[78]
port 246 nsew signal input
flabel metal2 s 405986 -960 406098 480 0 FreeSans 448 90 0 0 la_data_in[79]
port 247 nsew signal input
flabel metal2 s 150594 -960 150706 480 0 FreeSans 448 90 0 0 la_data_in[7]
port 248 nsew signal input
flabel metal2 s 409574 -960 409686 480 0 FreeSans 448 90 0 0 la_data_in[80]
port 249 nsew signal input
flabel metal2 s 413070 -960 413182 480 0 FreeSans 448 90 0 0 la_data_in[81]
port 250 nsew signal input
flabel metal2 s 416658 -960 416770 480 0 FreeSans 448 90 0 0 la_data_in[82]
port 251 nsew signal input
flabel metal2 s 420154 -960 420266 480 0 FreeSans 448 90 0 0 la_data_in[83]
port 252 nsew signal input
flabel metal2 s 423742 -960 423854 480 0 FreeSans 448 90 0 0 la_data_in[84]
port 253 nsew signal input
flabel metal2 s 427238 -960 427350 480 0 FreeSans 448 90 0 0 la_data_in[85]
port 254 nsew signal input
flabel metal2 s 430826 -960 430938 480 0 FreeSans 448 90 0 0 la_data_in[86]
port 255 nsew signal input
flabel metal2 s 434414 -960 434526 480 0 FreeSans 448 90 0 0 la_data_in[87]
port 256 nsew signal input
flabel metal2 s 437910 -960 438022 480 0 FreeSans 448 90 0 0 la_data_in[88]
port 257 nsew signal input
flabel metal2 s 441498 -960 441610 480 0 FreeSans 448 90 0 0 la_data_in[89]
port 258 nsew signal input
flabel metal2 s 154182 -960 154294 480 0 FreeSans 448 90 0 0 la_data_in[8]
port 259 nsew signal input
flabel metal2 s 444994 -960 445106 480 0 FreeSans 448 90 0 0 la_data_in[90]
port 260 nsew signal input
flabel metal2 s 448582 -960 448694 480 0 FreeSans 448 90 0 0 la_data_in[91]
port 261 nsew signal input
flabel metal2 s 452078 -960 452190 480 0 FreeSans 448 90 0 0 la_data_in[92]
port 262 nsew signal input
flabel metal2 s 455666 -960 455778 480 0 FreeSans 448 90 0 0 la_data_in[93]
port 263 nsew signal input
flabel metal2 s 459162 -960 459274 480 0 FreeSans 448 90 0 0 la_data_in[94]
port 264 nsew signal input
flabel metal2 s 462750 -960 462862 480 0 FreeSans 448 90 0 0 la_data_in[95]
port 265 nsew signal input
flabel metal2 s 466246 -960 466358 480 0 FreeSans 448 90 0 0 la_data_in[96]
port 266 nsew signal input
flabel metal2 s 469834 -960 469946 480 0 FreeSans 448 90 0 0 la_data_in[97]
port 267 nsew signal input
flabel metal2 s 473422 -960 473534 480 0 FreeSans 448 90 0 0 la_data_in[98]
port 268 nsew signal input
flabel metal2 s 476918 -960 477030 480 0 FreeSans 448 90 0 0 la_data_in[99]
port 269 nsew signal input
flabel metal2 s 157770 -960 157882 480 0 FreeSans 448 90 0 0 la_data_in[9]
port 270 nsew signal input
flabel metal2 s 126950 -960 127062 480 0 FreeSans 448 90 0 0 la_data_out[0]
port 271 nsew signal tristate
flabel metal2 s 481702 -960 481814 480 0 FreeSans 448 90 0 0 la_data_out[100]
port 272 nsew signal tristate
flabel metal2 s 485198 -960 485310 480 0 FreeSans 448 90 0 0 la_data_out[101]
port 273 nsew signal tristate
flabel metal2 s 488786 -960 488898 480 0 FreeSans 448 90 0 0 la_data_out[102]
port 274 nsew signal tristate
flabel metal2 s 492282 -960 492394 480 0 FreeSans 448 90 0 0 la_data_out[103]
port 275 nsew signal tristate
flabel metal2 s 495870 -960 495982 480 0 FreeSans 448 90 0 0 la_data_out[104]
port 276 nsew signal tristate
flabel metal2 s 499366 -960 499478 480 0 FreeSans 448 90 0 0 la_data_out[105]
port 277 nsew signal tristate
flabel metal2 s 502954 -960 503066 480 0 FreeSans 448 90 0 0 la_data_out[106]
port 278 nsew signal tristate
flabel metal2 s 506450 -960 506562 480 0 FreeSans 448 90 0 0 la_data_out[107]
port 279 nsew signal tristate
flabel metal2 s 510038 -960 510150 480 0 FreeSans 448 90 0 0 la_data_out[108]
port 280 nsew signal tristate
flabel metal2 s 513534 -960 513646 480 0 FreeSans 448 90 0 0 la_data_out[109]
port 281 nsew signal tristate
flabel metal2 s 162462 -960 162574 480 0 FreeSans 448 90 0 0 la_data_out[10]
port 282 nsew signal tristate
flabel metal2 s 517122 -960 517234 480 0 FreeSans 448 90 0 0 la_data_out[110]
port 283 nsew signal tristate
flabel metal2 s 520710 -960 520822 480 0 FreeSans 448 90 0 0 la_data_out[111]
port 284 nsew signal tristate
flabel metal2 s 524206 -960 524318 480 0 FreeSans 448 90 0 0 la_data_out[112]
port 285 nsew signal tristate
flabel metal2 s 527794 -960 527906 480 0 FreeSans 448 90 0 0 la_data_out[113]
port 286 nsew signal tristate
flabel metal2 s 531290 -960 531402 480 0 FreeSans 448 90 0 0 la_data_out[114]
port 287 nsew signal tristate
flabel metal2 s 534878 -960 534990 480 0 FreeSans 448 90 0 0 la_data_out[115]
port 288 nsew signal tristate
flabel metal2 s 538374 -960 538486 480 0 FreeSans 448 90 0 0 la_data_out[116]
port 289 nsew signal tristate
flabel metal2 s 541962 -960 542074 480 0 FreeSans 448 90 0 0 la_data_out[117]
port 290 nsew signal tristate
flabel metal2 s 545458 -960 545570 480 0 FreeSans 448 90 0 0 la_data_out[118]
port 291 nsew signal tristate
flabel metal2 s 549046 -960 549158 480 0 FreeSans 448 90 0 0 la_data_out[119]
port 292 nsew signal tristate
flabel metal2 s 166050 -960 166162 480 0 FreeSans 448 90 0 0 la_data_out[11]
port 293 nsew signal tristate
flabel metal2 s 552634 -960 552746 480 0 FreeSans 448 90 0 0 la_data_out[120]
port 294 nsew signal tristate
flabel metal2 s 556130 -960 556242 480 0 FreeSans 448 90 0 0 la_data_out[121]
port 295 nsew signal tristate
flabel metal2 s 559718 -960 559830 480 0 FreeSans 448 90 0 0 la_data_out[122]
port 296 nsew signal tristate
flabel metal2 s 563214 -960 563326 480 0 FreeSans 448 90 0 0 la_data_out[123]
port 297 nsew signal tristate
flabel metal2 s 566802 -960 566914 480 0 FreeSans 448 90 0 0 la_data_out[124]
port 298 nsew signal tristate
flabel metal2 s 570298 -960 570410 480 0 FreeSans 448 90 0 0 la_data_out[125]
port 299 nsew signal tristate
flabel metal2 s 573886 -960 573998 480 0 FreeSans 448 90 0 0 la_data_out[126]
port 300 nsew signal tristate
flabel metal2 s 577382 -960 577494 480 0 FreeSans 448 90 0 0 la_data_out[127]
port 301 nsew signal tristate
flabel metal2 s 169546 -960 169658 480 0 FreeSans 448 90 0 0 la_data_out[12]
port 302 nsew signal tristate
flabel metal2 s 173134 -960 173246 480 0 FreeSans 448 90 0 0 la_data_out[13]
port 303 nsew signal tristate
flabel metal2 s 176630 -960 176742 480 0 FreeSans 448 90 0 0 la_data_out[14]
port 304 nsew signal tristate
flabel metal2 s 180218 -960 180330 480 0 FreeSans 448 90 0 0 la_data_out[15]
port 305 nsew signal tristate
flabel metal2 s 183714 -960 183826 480 0 FreeSans 448 90 0 0 la_data_out[16]
port 306 nsew signal tristate
flabel metal2 s 187302 -960 187414 480 0 FreeSans 448 90 0 0 la_data_out[17]
port 307 nsew signal tristate
flabel metal2 s 190798 -960 190910 480 0 FreeSans 448 90 0 0 la_data_out[18]
port 308 nsew signal tristate
flabel metal2 s 194386 -960 194498 480 0 FreeSans 448 90 0 0 la_data_out[19]
port 309 nsew signal tristate
flabel metal2 s 130538 -960 130650 480 0 FreeSans 448 90 0 0 la_data_out[1]
port 310 nsew signal tristate
flabel metal2 s 197882 -960 197994 480 0 FreeSans 448 90 0 0 la_data_out[20]
port 311 nsew signal tristate
flabel metal2 s 201470 -960 201582 480 0 FreeSans 448 90 0 0 la_data_out[21]
port 312 nsew signal tristate
flabel metal2 s 205058 -960 205170 480 0 FreeSans 448 90 0 0 la_data_out[22]
port 313 nsew signal tristate
flabel metal2 s 208554 -960 208666 480 0 FreeSans 448 90 0 0 la_data_out[23]
port 314 nsew signal tristate
flabel metal2 s 212142 -960 212254 480 0 FreeSans 448 90 0 0 la_data_out[24]
port 315 nsew signal tristate
flabel metal2 s 215638 -960 215750 480 0 FreeSans 448 90 0 0 la_data_out[25]
port 316 nsew signal tristate
flabel metal2 s 219226 -960 219338 480 0 FreeSans 448 90 0 0 la_data_out[26]
port 317 nsew signal tristate
flabel metal2 s 222722 -960 222834 480 0 FreeSans 448 90 0 0 la_data_out[27]
port 318 nsew signal tristate
flabel metal2 s 226310 -960 226422 480 0 FreeSans 448 90 0 0 la_data_out[28]
port 319 nsew signal tristate
flabel metal2 s 229806 -960 229918 480 0 FreeSans 448 90 0 0 la_data_out[29]
port 320 nsew signal tristate
flabel metal2 s 134126 -960 134238 480 0 FreeSans 448 90 0 0 la_data_out[2]
port 321 nsew signal tristate
flabel metal2 s 233394 -960 233506 480 0 FreeSans 448 90 0 0 la_data_out[30]
port 322 nsew signal tristate
flabel metal2 s 236982 -960 237094 480 0 FreeSans 448 90 0 0 la_data_out[31]
port 323 nsew signal tristate
flabel metal2 s 240478 -960 240590 480 0 FreeSans 448 90 0 0 la_data_out[32]
port 324 nsew signal tristate
flabel metal2 s 244066 -960 244178 480 0 FreeSans 448 90 0 0 la_data_out[33]
port 325 nsew signal tristate
flabel metal2 s 247562 -960 247674 480 0 FreeSans 448 90 0 0 la_data_out[34]
port 326 nsew signal tristate
flabel metal2 s 251150 -960 251262 480 0 FreeSans 448 90 0 0 la_data_out[35]
port 327 nsew signal tristate
flabel metal2 s 254646 -960 254758 480 0 FreeSans 448 90 0 0 la_data_out[36]
port 328 nsew signal tristate
flabel metal2 s 258234 -960 258346 480 0 FreeSans 448 90 0 0 la_data_out[37]
port 329 nsew signal tristate
flabel metal2 s 261730 -960 261842 480 0 FreeSans 448 90 0 0 la_data_out[38]
port 330 nsew signal tristate
flabel metal2 s 265318 -960 265430 480 0 FreeSans 448 90 0 0 la_data_out[39]
port 331 nsew signal tristate
flabel metal2 s 137622 -960 137734 480 0 FreeSans 448 90 0 0 la_data_out[3]
port 332 nsew signal tristate
flabel metal2 s 268814 -960 268926 480 0 FreeSans 448 90 0 0 la_data_out[40]
port 333 nsew signal tristate
flabel metal2 s 272402 -960 272514 480 0 FreeSans 448 90 0 0 la_data_out[41]
port 334 nsew signal tristate
flabel metal2 s 275990 -960 276102 480 0 FreeSans 448 90 0 0 la_data_out[42]
port 335 nsew signal tristate
flabel metal2 s 279486 -960 279598 480 0 FreeSans 448 90 0 0 la_data_out[43]
port 336 nsew signal tristate
flabel metal2 s 283074 -960 283186 480 0 FreeSans 448 90 0 0 la_data_out[44]
port 337 nsew signal tristate
flabel metal2 s 286570 -960 286682 480 0 FreeSans 448 90 0 0 la_data_out[45]
port 338 nsew signal tristate
flabel metal2 s 290158 -960 290270 480 0 FreeSans 448 90 0 0 la_data_out[46]
port 339 nsew signal tristate
flabel metal2 s 293654 -960 293766 480 0 FreeSans 448 90 0 0 la_data_out[47]
port 340 nsew signal tristate
flabel metal2 s 297242 -960 297354 480 0 FreeSans 448 90 0 0 la_data_out[48]
port 341 nsew signal tristate
flabel metal2 s 300738 -960 300850 480 0 FreeSans 448 90 0 0 la_data_out[49]
port 342 nsew signal tristate
flabel metal2 s 141210 -960 141322 480 0 FreeSans 448 90 0 0 la_data_out[4]
port 343 nsew signal tristate
flabel metal2 s 304326 -960 304438 480 0 FreeSans 448 90 0 0 la_data_out[50]
port 344 nsew signal tristate
flabel metal2 s 307914 -960 308026 480 0 FreeSans 448 90 0 0 la_data_out[51]
port 345 nsew signal tristate
flabel metal2 s 311410 -960 311522 480 0 FreeSans 448 90 0 0 la_data_out[52]
port 346 nsew signal tristate
flabel metal2 s 314998 -960 315110 480 0 FreeSans 448 90 0 0 la_data_out[53]
port 347 nsew signal tristate
flabel metal2 s 318494 -960 318606 480 0 FreeSans 448 90 0 0 la_data_out[54]
port 348 nsew signal tristate
flabel metal2 s 322082 -960 322194 480 0 FreeSans 448 90 0 0 la_data_out[55]
port 349 nsew signal tristate
flabel metal2 s 325578 -960 325690 480 0 FreeSans 448 90 0 0 la_data_out[56]
port 350 nsew signal tristate
flabel metal2 s 329166 -960 329278 480 0 FreeSans 448 90 0 0 la_data_out[57]
port 351 nsew signal tristate
flabel metal2 s 332662 -960 332774 480 0 FreeSans 448 90 0 0 la_data_out[58]
port 352 nsew signal tristate
flabel metal2 s 336250 -960 336362 480 0 FreeSans 448 90 0 0 la_data_out[59]
port 353 nsew signal tristate
flabel metal2 s 144706 -960 144818 480 0 FreeSans 448 90 0 0 la_data_out[5]
port 354 nsew signal tristate
flabel metal2 s 339838 -960 339950 480 0 FreeSans 448 90 0 0 la_data_out[60]
port 355 nsew signal tristate
flabel metal2 s 343334 -960 343446 480 0 FreeSans 448 90 0 0 la_data_out[61]
port 356 nsew signal tristate
flabel metal2 s 346922 -960 347034 480 0 FreeSans 448 90 0 0 la_data_out[62]
port 357 nsew signal tristate
flabel metal2 s 350418 -960 350530 480 0 FreeSans 448 90 0 0 la_data_out[63]
port 358 nsew signal tristate
flabel metal2 s 354006 -960 354118 480 0 FreeSans 448 90 0 0 la_data_out[64]
port 359 nsew signal tristate
flabel metal2 s 357502 -960 357614 480 0 FreeSans 448 90 0 0 la_data_out[65]
port 360 nsew signal tristate
flabel metal2 s 361090 -960 361202 480 0 FreeSans 448 90 0 0 la_data_out[66]
port 361 nsew signal tristate
flabel metal2 s 364586 -960 364698 480 0 FreeSans 448 90 0 0 la_data_out[67]
port 362 nsew signal tristate
flabel metal2 s 368174 -960 368286 480 0 FreeSans 448 90 0 0 la_data_out[68]
port 363 nsew signal tristate
flabel metal2 s 371670 -960 371782 480 0 FreeSans 448 90 0 0 la_data_out[69]
port 364 nsew signal tristate
flabel metal2 s 148294 -960 148406 480 0 FreeSans 448 90 0 0 la_data_out[6]
port 365 nsew signal tristate
flabel metal2 s 375258 -960 375370 480 0 FreeSans 448 90 0 0 la_data_out[70]
port 366 nsew signal tristate
flabel metal2 s 378846 -960 378958 480 0 FreeSans 448 90 0 0 la_data_out[71]
port 367 nsew signal tristate
flabel metal2 s 382342 -960 382454 480 0 FreeSans 448 90 0 0 la_data_out[72]
port 368 nsew signal tristate
flabel metal2 s 385930 -960 386042 480 0 FreeSans 448 90 0 0 la_data_out[73]
port 369 nsew signal tristate
flabel metal2 s 389426 -960 389538 480 0 FreeSans 448 90 0 0 la_data_out[74]
port 370 nsew signal tristate
flabel metal2 s 393014 -960 393126 480 0 FreeSans 448 90 0 0 la_data_out[75]
port 371 nsew signal tristate
flabel metal2 s 396510 -960 396622 480 0 FreeSans 448 90 0 0 la_data_out[76]
port 372 nsew signal tristate
flabel metal2 s 400098 -960 400210 480 0 FreeSans 448 90 0 0 la_data_out[77]
port 373 nsew signal tristate
flabel metal2 s 403594 -960 403706 480 0 FreeSans 448 90 0 0 la_data_out[78]
port 374 nsew signal tristate
flabel metal2 s 407182 -960 407294 480 0 FreeSans 448 90 0 0 la_data_out[79]
port 375 nsew signal tristate
flabel metal2 s 151790 -960 151902 480 0 FreeSans 448 90 0 0 la_data_out[7]
port 376 nsew signal tristate
flabel metal2 s 410770 -960 410882 480 0 FreeSans 448 90 0 0 la_data_out[80]
port 377 nsew signal tristate
flabel metal2 s 414266 -960 414378 480 0 FreeSans 448 90 0 0 la_data_out[81]
port 378 nsew signal tristate
flabel metal2 s 417854 -960 417966 480 0 FreeSans 448 90 0 0 la_data_out[82]
port 379 nsew signal tristate
flabel metal2 s 421350 -960 421462 480 0 FreeSans 448 90 0 0 la_data_out[83]
port 380 nsew signal tristate
flabel metal2 s 424938 -960 425050 480 0 FreeSans 448 90 0 0 la_data_out[84]
port 381 nsew signal tristate
flabel metal2 s 428434 -960 428546 480 0 FreeSans 448 90 0 0 la_data_out[85]
port 382 nsew signal tristate
flabel metal2 s 432022 -960 432134 480 0 FreeSans 448 90 0 0 la_data_out[86]
port 383 nsew signal tristate
flabel metal2 s 435518 -960 435630 480 0 FreeSans 448 90 0 0 la_data_out[87]
port 384 nsew signal tristate
flabel metal2 s 439106 -960 439218 480 0 FreeSans 448 90 0 0 la_data_out[88]
port 385 nsew signal tristate
flabel metal2 s 442602 -960 442714 480 0 FreeSans 448 90 0 0 la_data_out[89]
port 386 nsew signal tristate
flabel metal2 s 155378 -960 155490 480 0 FreeSans 448 90 0 0 la_data_out[8]
port 387 nsew signal tristate
flabel metal2 s 446190 -960 446302 480 0 FreeSans 448 90 0 0 la_data_out[90]
port 388 nsew signal tristate
flabel metal2 s 449778 -960 449890 480 0 FreeSans 448 90 0 0 la_data_out[91]
port 389 nsew signal tristate
flabel metal2 s 453274 -960 453386 480 0 FreeSans 448 90 0 0 la_data_out[92]
port 390 nsew signal tristate
flabel metal2 s 456862 -960 456974 480 0 FreeSans 448 90 0 0 la_data_out[93]
port 391 nsew signal tristate
flabel metal2 s 460358 -960 460470 480 0 FreeSans 448 90 0 0 la_data_out[94]
port 392 nsew signal tristate
flabel metal2 s 463946 -960 464058 480 0 FreeSans 448 90 0 0 la_data_out[95]
port 393 nsew signal tristate
flabel metal2 s 467442 -960 467554 480 0 FreeSans 448 90 0 0 la_data_out[96]
port 394 nsew signal tristate
flabel metal2 s 471030 -960 471142 480 0 FreeSans 448 90 0 0 la_data_out[97]
port 395 nsew signal tristate
flabel metal2 s 474526 -960 474638 480 0 FreeSans 448 90 0 0 la_data_out[98]
port 396 nsew signal tristate
flabel metal2 s 478114 -960 478226 480 0 FreeSans 448 90 0 0 la_data_out[99]
port 397 nsew signal tristate
flabel metal2 s 158874 -960 158986 480 0 FreeSans 448 90 0 0 la_data_out[9]
port 398 nsew signal tristate
flabel metal2 s 128146 -960 128258 480 0 FreeSans 448 90 0 0 la_oenb[0]
port 399 nsew signal input
flabel metal2 s 482806 -960 482918 480 0 FreeSans 448 90 0 0 la_oenb[100]
port 400 nsew signal input
flabel metal2 s 486394 -960 486506 480 0 FreeSans 448 90 0 0 la_oenb[101]
port 401 nsew signal input
flabel metal2 s 489890 -960 490002 480 0 FreeSans 448 90 0 0 la_oenb[102]
port 402 nsew signal input
flabel metal2 s 493478 -960 493590 480 0 FreeSans 448 90 0 0 la_oenb[103]
port 403 nsew signal input
flabel metal2 s 497066 -960 497178 480 0 FreeSans 448 90 0 0 la_oenb[104]
port 404 nsew signal input
flabel metal2 s 500562 -960 500674 480 0 FreeSans 448 90 0 0 la_oenb[105]
port 405 nsew signal input
flabel metal2 s 504150 -960 504262 480 0 FreeSans 448 90 0 0 la_oenb[106]
port 406 nsew signal input
flabel metal2 s 507646 -960 507758 480 0 FreeSans 448 90 0 0 la_oenb[107]
port 407 nsew signal input
flabel metal2 s 511234 -960 511346 480 0 FreeSans 448 90 0 0 la_oenb[108]
port 408 nsew signal input
flabel metal2 s 514730 -960 514842 480 0 FreeSans 448 90 0 0 la_oenb[109]
port 409 nsew signal input
flabel metal2 s 163658 -960 163770 480 0 FreeSans 448 90 0 0 la_oenb[10]
port 410 nsew signal input
flabel metal2 s 518318 -960 518430 480 0 FreeSans 448 90 0 0 la_oenb[110]
port 411 nsew signal input
flabel metal2 s 521814 -960 521926 480 0 FreeSans 448 90 0 0 la_oenb[111]
port 412 nsew signal input
flabel metal2 s 525402 -960 525514 480 0 FreeSans 448 90 0 0 la_oenb[112]
port 413 nsew signal input
flabel metal2 s 528990 -960 529102 480 0 FreeSans 448 90 0 0 la_oenb[113]
port 414 nsew signal input
flabel metal2 s 532486 -960 532598 480 0 FreeSans 448 90 0 0 la_oenb[114]
port 415 nsew signal input
flabel metal2 s 536074 -960 536186 480 0 FreeSans 448 90 0 0 la_oenb[115]
port 416 nsew signal input
flabel metal2 s 539570 -960 539682 480 0 FreeSans 448 90 0 0 la_oenb[116]
port 417 nsew signal input
flabel metal2 s 543158 -960 543270 480 0 FreeSans 448 90 0 0 la_oenb[117]
port 418 nsew signal input
flabel metal2 s 546654 -960 546766 480 0 FreeSans 448 90 0 0 la_oenb[118]
port 419 nsew signal input
flabel metal2 s 550242 -960 550354 480 0 FreeSans 448 90 0 0 la_oenb[119]
port 420 nsew signal input
flabel metal2 s 167154 -960 167266 480 0 FreeSans 448 90 0 0 la_oenb[11]
port 421 nsew signal input
flabel metal2 s 553738 -960 553850 480 0 FreeSans 448 90 0 0 la_oenb[120]
port 422 nsew signal input
flabel metal2 s 557326 -960 557438 480 0 FreeSans 448 90 0 0 la_oenb[121]
port 423 nsew signal input
flabel metal2 s 560822 -960 560934 480 0 FreeSans 448 90 0 0 la_oenb[122]
port 424 nsew signal input
flabel metal2 s 564410 -960 564522 480 0 FreeSans 448 90 0 0 la_oenb[123]
port 425 nsew signal input
flabel metal2 s 567998 -960 568110 480 0 FreeSans 448 90 0 0 la_oenb[124]
port 426 nsew signal input
flabel metal2 s 571494 -960 571606 480 0 FreeSans 448 90 0 0 la_oenb[125]
port 427 nsew signal input
flabel metal2 s 575082 -960 575194 480 0 FreeSans 448 90 0 0 la_oenb[126]
port 428 nsew signal input
flabel metal2 s 578578 -960 578690 480 0 FreeSans 448 90 0 0 la_oenb[127]
port 429 nsew signal input
flabel metal2 s 170742 -960 170854 480 0 FreeSans 448 90 0 0 la_oenb[12]
port 430 nsew signal input
flabel metal2 s 174238 -960 174350 480 0 FreeSans 448 90 0 0 la_oenb[13]
port 431 nsew signal input
flabel metal2 s 177826 -960 177938 480 0 FreeSans 448 90 0 0 la_oenb[14]
port 432 nsew signal input
flabel metal2 s 181414 -960 181526 480 0 FreeSans 448 90 0 0 la_oenb[15]
port 433 nsew signal input
flabel metal2 s 184910 -960 185022 480 0 FreeSans 448 90 0 0 la_oenb[16]
port 434 nsew signal input
flabel metal2 s 188498 -960 188610 480 0 FreeSans 448 90 0 0 la_oenb[17]
port 435 nsew signal input
flabel metal2 s 191994 -960 192106 480 0 FreeSans 448 90 0 0 la_oenb[18]
port 436 nsew signal input
flabel metal2 s 195582 -960 195694 480 0 FreeSans 448 90 0 0 la_oenb[19]
port 437 nsew signal input
flabel metal2 s 131734 -960 131846 480 0 FreeSans 448 90 0 0 la_oenb[1]
port 438 nsew signal input
flabel metal2 s 199078 -960 199190 480 0 FreeSans 448 90 0 0 la_oenb[20]
port 439 nsew signal input
flabel metal2 s 202666 -960 202778 480 0 FreeSans 448 90 0 0 la_oenb[21]
port 440 nsew signal input
flabel metal2 s 206162 -960 206274 480 0 FreeSans 448 90 0 0 la_oenb[22]
port 441 nsew signal input
flabel metal2 s 209750 -960 209862 480 0 FreeSans 448 90 0 0 la_oenb[23]
port 442 nsew signal input
flabel metal2 s 213338 -960 213450 480 0 FreeSans 448 90 0 0 la_oenb[24]
port 443 nsew signal input
flabel metal2 s 216834 -960 216946 480 0 FreeSans 448 90 0 0 la_oenb[25]
port 444 nsew signal input
flabel metal2 s 220422 -960 220534 480 0 FreeSans 448 90 0 0 la_oenb[26]
port 445 nsew signal input
flabel metal2 s 223918 -960 224030 480 0 FreeSans 448 90 0 0 la_oenb[27]
port 446 nsew signal input
flabel metal2 s 227506 -960 227618 480 0 FreeSans 448 90 0 0 la_oenb[28]
port 447 nsew signal input
flabel metal2 s 231002 -960 231114 480 0 FreeSans 448 90 0 0 la_oenb[29]
port 448 nsew signal input
flabel metal2 s 135230 -960 135342 480 0 FreeSans 448 90 0 0 la_oenb[2]
port 449 nsew signal input
flabel metal2 s 234590 -960 234702 480 0 FreeSans 448 90 0 0 la_oenb[30]
port 450 nsew signal input
flabel metal2 s 238086 -960 238198 480 0 FreeSans 448 90 0 0 la_oenb[31]
port 451 nsew signal input
flabel metal2 s 241674 -960 241786 480 0 FreeSans 448 90 0 0 la_oenb[32]
port 452 nsew signal input
flabel metal2 s 245170 -960 245282 480 0 FreeSans 448 90 0 0 la_oenb[33]
port 453 nsew signal input
flabel metal2 s 248758 -960 248870 480 0 FreeSans 448 90 0 0 la_oenb[34]
port 454 nsew signal input
flabel metal2 s 252346 -960 252458 480 0 FreeSans 448 90 0 0 la_oenb[35]
port 455 nsew signal input
flabel metal2 s 255842 -960 255954 480 0 FreeSans 448 90 0 0 la_oenb[36]
port 456 nsew signal input
flabel metal2 s 259430 -960 259542 480 0 FreeSans 448 90 0 0 la_oenb[37]
port 457 nsew signal input
flabel metal2 s 262926 -960 263038 480 0 FreeSans 448 90 0 0 la_oenb[38]
port 458 nsew signal input
flabel metal2 s 266514 -960 266626 480 0 FreeSans 448 90 0 0 la_oenb[39]
port 459 nsew signal input
flabel metal2 s 138818 -960 138930 480 0 FreeSans 448 90 0 0 la_oenb[3]
port 460 nsew signal input
flabel metal2 s 270010 -960 270122 480 0 FreeSans 448 90 0 0 la_oenb[40]
port 461 nsew signal input
flabel metal2 s 273598 -960 273710 480 0 FreeSans 448 90 0 0 la_oenb[41]
port 462 nsew signal input
flabel metal2 s 277094 -960 277206 480 0 FreeSans 448 90 0 0 la_oenb[42]
port 463 nsew signal input
flabel metal2 s 280682 -960 280794 480 0 FreeSans 448 90 0 0 la_oenb[43]
port 464 nsew signal input
flabel metal2 s 284270 -960 284382 480 0 FreeSans 448 90 0 0 la_oenb[44]
port 465 nsew signal input
flabel metal2 s 287766 -960 287878 480 0 FreeSans 448 90 0 0 la_oenb[45]
port 466 nsew signal input
flabel metal2 s 291354 -960 291466 480 0 FreeSans 448 90 0 0 la_oenb[46]
port 467 nsew signal input
flabel metal2 s 294850 -960 294962 480 0 FreeSans 448 90 0 0 la_oenb[47]
port 468 nsew signal input
flabel metal2 s 298438 -960 298550 480 0 FreeSans 448 90 0 0 la_oenb[48]
port 469 nsew signal input
flabel metal2 s 301934 -960 302046 480 0 FreeSans 448 90 0 0 la_oenb[49]
port 470 nsew signal input
flabel metal2 s 142406 -960 142518 480 0 FreeSans 448 90 0 0 la_oenb[4]
port 471 nsew signal input
flabel metal2 s 305522 -960 305634 480 0 FreeSans 448 90 0 0 la_oenb[50]
port 472 nsew signal input
flabel metal2 s 309018 -960 309130 480 0 FreeSans 448 90 0 0 la_oenb[51]
port 473 nsew signal input
flabel metal2 s 312606 -960 312718 480 0 FreeSans 448 90 0 0 la_oenb[52]
port 474 nsew signal input
flabel metal2 s 316194 -960 316306 480 0 FreeSans 448 90 0 0 la_oenb[53]
port 475 nsew signal input
flabel metal2 s 319690 -960 319802 480 0 FreeSans 448 90 0 0 la_oenb[54]
port 476 nsew signal input
flabel metal2 s 323278 -960 323390 480 0 FreeSans 448 90 0 0 la_oenb[55]
port 477 nsew signal input
flabel metal2 s 326774 -960 326886 480 0 FreeSans 448 90 0 0 la_oenb[56]
port 478 nsew signal input
flabel metal2 s 330362 -960 330474 480 0 FreeSans 448 90 0 0 la_oenb[57]
port 479 nsew signal input
flabel metal2 s 333858 -960 333970 480 0 FreeSans 448 90 0 0 la_oenb[58]
port 480 nsew signal input
flabel metal2 s 337446 -960 337558 480 0 FreeSans 448 90 0 0 la_oenb[59]
port 481 nsew signal input
flabel metal2 s 145902 -960 146014 480 0 FreeSans 448 90 0 0 la_oenb[5]
port 482 nsew signal input
flabel metal2 s 340942 -960 341054 480 0 FreeSans 448 90 0 0 la_oenb[60]
port 483 nsew signal input
flabel metal2 s 344530 -960 344642 480 0 FreeSans 448 90 0 0 la_oenb[61]
port 484 nsew signal input
flabel metal2 s 348026 -960 348138 480 0 FreeSans 448 90 0 0 la_oenb[62]
port 485 nsew signal input
flabel metal2 s 351614 -960 351726 480 0 FreeSans 448 90 0 0 la_oenb[63]
port 486 nsew signal input
flabel metal2 s 355202 -960 355314 480 0 FreeSans 448 90 0 0 la_oenb[64]
port 487 nsew signal input
flabel metal2 s 358698 -960 358810 480 0 FreeSans 448 90 0 0 la_oenb[65]
port 488 nsew signal input
flabel metal2 s 362286 -960 362398 480 0 FreeSans 448 90 0 0 la_oenb[66]
port 489 nsew signal input
flabel metal2 s 365782 -960 365894 480 0 FreeSans 448 90 0 0 la_oenb[67]
port 490 nsew signal input
flabel metal2 s 369370 -960 369482 480 0 FreeSans 448 90 0 0 la_oenb[68]
port 491 nsew signal input
flabel metal2 s 372866 -960 372978 480 0 FreeSans 448 90 0 0 la_oenb[69]
port 492 nsew signal input
flabel metal2 s 149490 -960 149602 480 0 FreeSans 448 90 0 0 la_oenb[6]
port 493 nsew signal input
flabel metal2 s 376454 -960 376566 480 0 FreeSans 448 90 0 0 la_oenb[70]
port 494 nsew signal input
flabel metal2 s 379950 -960 380062 480 0 FreeSans 448 90 0 0 la_oenb[71]
port 495 nsew signal input
flabel metal2 s 383538 -960 383650 480 0 FreeSans 448 90 0 0 la_oenb[72]
port 496 nsew signal input
flabel metal2 s 387126 -960 387238 480 0 FreeSans 448 90 0 0 la_oenb[73]
port 497 nsew signal input
flabel metal2 s 390622 -960 390734 480 0 FreeSans 448 90 0 0 la_oenb[74]
port 498 nsew signal input
flabel metal2 s 394210 -960 394322 480 0 FreeSans 448 90 0 0 la_oenb[75]
port 499 nsew signal input
flabel metal2 s 397706 -960 397818 480 0 FreeSans 448 90 0 0 la_oenb[76]
port 500 nsew signal input
flabel metal2 s 401294 -960 401406 480 0 FreeSans 448 90 0 0 la_oenb[77]
port 501 nsew signal input
flabel metal2 s 404790 -960 404902 480 0 FreeSans 448 90 0 0 la_oenb[78]
port 502 nsew signal input
flabel metal2 s 408378 -960 408490 480 0 FreeSans 448 90 0 0 la_oenb[79]
port 503 nsew signal input
flabel metal2 s 152986 -960 153098 480 0 FreeSans 448 90 0 0 la_oenb[7]
port 504 nsew signal input
flabel metal2 s 411874 -960 411986 480 0 FreeSans 448 90 0 0 la_oenb[80]
port 505 nsew signal input
flabel metal2 s 415462 -960 415574 480 0 FreeSans 448 90 0 0 la_oenb[81]
port 506 nsew signal input
flabel metal2 s 418958 -960 419070 480 0 FreeSans 448 90 0 0 la_oenb[82]
port 507 nsew signal input
flabel metal2 s 422546 -960 422658 480 0 FreeSans 448 90 0 0 la_oenb[83]
port 508 nsew signal input
flabel metal2 s 426134 -960 426246 480 0 FreeSans 448 90 0 0 la_oenb[84]
port 509 nsew signal input
flabel metal2 s 429630 -960 429742 480 0 FreeSans 448 90 0 0 la_oenb[85]
port 510 nsew signal input
flabel metal2 s 433218 -960 433330 480 0 FreeSans 448 90 0 0 la_oenb[86]
port 511 nsew signal input
flabel metal2 s 436714 -960 436826 480 0 FreeSans 448 90 0 0 la_oenb[87]
port 512 nsew signal input
flabel metal2 s 440302 -960 440414 480 0 FreeSans 448 90 0 0 la_oenb[88]
port 513 nsew signal input
flabel metal2 s 443798 -960 443910 480 0 FreeSans 448 90 0 0 la_oenb[89]
port 514 nsew signal input
flabel metal2 s 156574 -960 156686 480 0 FreeSans 448 90 0 0 la_oenb[8]
port 515 nsew signal input
flabel metal2 s 447386 -960 447498 480 0 FreeSans 448 90 0 0 la_oenb[90]
port 516 nsew signal input
flabel metal2 s 450882 -960 450994 480 0 FreeSans 448 90 0 0 la_oenb[91]
port 517 nsew signal input
flabel metal2 s 454470 -960 454582 480 0 FreeSans 448 90 0 0 la_oenb[92]
port 518 nsew signal input
flabel metal2 s 458058 -960 458170 480 0 FreeSans 448 90 0 0 la_oenb[93]
port 519 nsew signal input
flabel metal2 s 461554 -960 461666 480 0 FreeSans 448 90 0 0 la_oenb[94]
port 520 nsew signal input
flabel metal2 s 465142 -960 465254 480 0 FreeSans 448 90 0 0 la_oenb[95]
port 521 nsew signal input
flabel metal2 s 468638 -960 468750 480 0 FreeSans 448 90 0 0 la_oenb[96]
port 522 nsew signal input
flabel metal2 s 472226 -960 472338 480 0 FreeSans 448 90 0 0 la_oenb[97]
port 523 nsew signal input
flabel metal2 s 475722 -960 475834 480 0 FreeSans 448 90 0 0 la_oenb[98]
port 524 nsew signal input
flabel metal2 s 479310 -960 479422 480 0 FreeSans 448 90 0 0 la_oenb[99]
port 525 nsew signal input
flabel metal2 s 160070 -960 160182 480 0 FreeSans 448 90 0 0 la_oenb[9]
port 526 nsew signal input
flabel metal2 s 579774 -960 579886 480 0 FreeSans 448 90 0 0 user_clock2
port 527 nsew signal input
flabel metal2 s 580970 -960 581082 480 0 FreeSans 448 90 0 0 user_irq[0]
port 528 nsew signal tristate
flabel metal2 s 582166 -960 582278 480 0 FreeSans 448 90 0 0 user_irq[1]
port 529 nsew signal tristate
flabel metal2 s 583362 -960 583474 480 0 FreeSans 448 90 0 0 user_irq[2]
port 530 nsew signal tristate
flabel metal4 s -2006 -934 -1386 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 -934 585930 -314 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 704250 585930 704870 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 585310 -934 585930 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 11866 592650 12486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 47866 592650 48486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 83866 592650 84486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 119866 592650 120486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 155866 592650 156486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 191866 592650 192486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 227866 592650 228486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 263866 592650 264486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 299866 592650 300486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 335866 592650 336486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 371866 592650 372486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 407866 592650 408486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 443866 592650 444486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 479866 592650 480486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 515866 592650 516486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 551866 592650 552486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 587866 592650 588486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 623866 592650 624486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 659866 592650 660486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 695866 592650 696486 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s -3926 -2854 -3306 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 -2854 587850 -2234 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 706170 587850 706790 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 587230 -2854 587850 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s -5846 -4774 -5226 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 -4774 589770 -4154 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 708090 589770 708710 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 589150 -4774 589770 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s -7766 -6694 -7146 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 -6694 591690 -6074 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 710010 591690 710630 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 591070 -6694 591690 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s -6806 -5734 -6186 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 -5734 590730 -5114 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 709050 590730 709670 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 590110 -5734 590730 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s -8726 -7654 -8106 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 -7654 592650 -7034 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 710970 592650 711590 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 592030 -7654 592650 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s -2966 -1894 -2346 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 -1894 586890 -1274 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 705210 586890 705830 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 586270 -1894 586890 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 582294 -7654 582914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 16366 592650 16986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 52366 592650 52986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 88366 592650 88986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 124366 592650 124986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 160366 592650 160986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 196366 592650 196986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 232366 592650 232986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 268366 592650 268986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 304366 592650 304986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 340366 592650 340986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 376366 592650 376986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 412366 592650 412986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 448366 592650 448986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 484366 592650 484986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 520366 592650 520986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 556366 592650 556986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 592366 592650 592986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 628366 592650 628986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 664366 592650 664986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 700366 592650 700986 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s -4886 -3814 -4266 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 -3814 588810 -3194 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 707130 588810 707750 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 588190 -3814 588810 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal2 s 542 -960 654 480 0 FreeSans 448 90 0 0 wb_clk_i
port 539 nsew signal input
flabel metal2 s 1646 -960 1758 480 0 FreeSans 448 90 0 0 wb_rst_i
port 540 nsew signal input
flabel metal2 s 2842 -960 2954 480 0 FreeSans 448 90 0 0 wbs_ack_o
port 541 nsew signal tristate
flabel metal2 s 7626 -960 7738 480 0 FreeSans 448 90 0 0 wbs_adr_i[0]
port 542 nsew signal input
flabel metal2 s 47830 -960 47942 480 0 FreeSans 448 90 0 0 wbs_adr_i[10]
port 543 nsew signal input
flabel metal2 s 51326 -960 51438 480 0 FreeSans 448 90 0 0 wbs_adr_i[11]
port 544 nsew signal input
flabel metal2 s 54914 -960 55026 480 0 FreeSans 448 90 0 0 wbs_adr_i[12]
port 545 nsew signal input
flabel metal2 s 58410 -960 58522 480 0 FreeSans 448 90 0 0 wbs_adr_i[13]
port 546 nsew signal input
flabel metal2 s 61998 -960 62110 480 0 FreeSans 448 90 0 0 wbs_adr_i[14]
port 547 nsew signal input
flabel metal2 s 65494 -960 65606 480 0 FreeSans 448 90 0 0 wbs_adr_i[15]
port 548 nsew signal input
flabel metal2 s 69082 -960 69194 480 0 FreeSans 448 90 0 0 wbs_adr_i[16]
port 549 nsew signal input
flabel metal2 s 72578 -960 72690 480 0 FreeSans 448 90 0 0 wbs_adr_i[17]
port 550 nsew signal input
flabel metal2 s 76166 -960 76278 480 0 FreeSans 448 90 0 0 wbs_adr_i[18]
port 551 nsew signal input
flabel metal2 s 79662 -960 79774 480 0 FreeSans 448 90 0 0 wbs_adr_i[19]
port 552 nsew signal input
flabel metal2 s 12318 -960 12430 480 0 FreeSans 448 90 0 0 wbs_adr_i[1]
port 553 nsew signal input
flabel metal2 s 83250 -960 83362 480 0 FreeSans 448 90 0 0 wbs_adr_i[20]
port 554 nsew signal input
flabel metal2 s 86838 -960 86950 480 0 FreeSans 448 90 0 0 wbs_adr_i[21]
port 555 nsew signal input
flabel metal2 s 90334 -960 90446 480 0 FreeSans 448 90 0 0 wbs_adr_i[22]
port 556 nsew signal input
flabel metal2 s 93922 -960 94034 480 0 FreeSans 448 90 0 0 wbs_adr_i[23]
port 557 nsew signal input
flabel metal2 s 97418 -960 97530 480 0 FreeSans 448 90 0 0 wbs_adr_i[24]
port 558 nsew signal input
flabel metal2 s 101006 -960 101118 480 0 FreeSans 448 90 0 0 wbs_adr_i[25]
port 559 nsew signal input
flabel metal2 s 104502 -960 104614 480 0 FreeSans 448 90 0 0 wbs_adr_i[26]
port 560 nsew signal input
flabel metal2 s 108090 -960 108202 480 0 FreeSans 448 90 0 0 wbs_adr_i[27]
port 561 nsew signal input
flabel metal2 s 111586 -960 111698 480 0 FreeSans 448 90 0 0 wbs_adr_i[28]
port 562 nsew signal input
flabel metal2 s 115174 -960 115286 480 0 FreeSans 448 90 0 0 wbs_adr_i[29]
port 563 nsew signal input
flabel metal2 s 17010 -960 17122 480 0 FreeSans 448 90 0 0 wbs_adr_i[2]
port 564 nsew signal input
flabel metal2 s 118762 -960 118874 480 0 FreeSans 448 90 0 0 wbs_adr_i[30]
port 565 nsew signal input
flabel metal2 s 122258 -960 122370 480 0 FreeSans 448 90 0 0 wbs_adr_i[31]
port 566 nsew signal input
flabel metal2 s 21794 -960 21906 480 0 FreeSans 448 90 0 0 wbs_adr_i[3]
port 567 nsew signal input
flabel metal2 s 26486 -960 26598 480 0 FreeSans 448 90 0 0 wbs_adr_i[4]
port 568 nsew signal input
flabel metal2 s 30074 -960 30186 480 0 FreeSans 448 90 0 0 wbs_adr_i[5]
port 569 nsew signal input
flabel metal2 s 33570 -960 33682 480 0 FreeSans 448 90 0 0 wbs_adr_i[6]
port 570 nsew signal input
flabel metal2 s 37158 -960 37270 480 0 FreeSans 448 90 0 0 wbs_adr_i[7]
port 571 nsew signal input
flabel metal2 s 40654 -960 40766 480 0 FreeSans 448 90 0 0 wbs_adr_i[8]
port 572 nsew signal input
flabel metal2 s 44242 -960 44354 480 0 FreeSans 448 90 0 0 wbs_adr_i[9]
port 573 nsew signal input
flabel metal2 s 4038 -960 4150 480 0 FreeSans 448 90 0 0 wbs_cyc_i
port 574 nsew signal input
flabel metal2 s 8730 -960 8842 480 0 FreeSans 448 90 0 0 wbs_dat_i[0]
port 575 nsew signal input
flabel metal2 s 48934 -960 49046 480 0 FreeSans 448 90 0 0 wbs_dat_i[10]
port 576 nsew signal input
flabel metal2 s 52522 -960 52634 480 0 FreeSans 448 90 0 0 wbs_dat_i[11]
port 577 nsew signal input
flabel metal2 s 56018 -960 56130 480 0 FreeSans 448 90 0 0 wbs_dat_i[12]
port 578 nsew signal input
flabel metal2 s 59606 -960 59718 480 0 FreeSans 448 90 0 0 wbs_dat_i[13]
port 579 nsew signal input
flabel metal2 s 63194 -960 63306 480 0 FreeSans 448 90 0 0 wbs_dat_i[14]
port 580 nsew signal input
flabel metal2 s 66690 -960 66802 480 0 FreeSans 448 90 0 0 wbs_dat_i[15]
port 581 nsew signal input
flabel metal2 s 70278 -960 70390 480 0 FreeSans 448 90 0 0 wbs_dat_i[16]
port 582 nsew signal input
flabel metal2 s 73774 -960 73886 480 0 FreeSans 448 90 0 0 wbs_dat_i[17]
port 583 nsew signal input
flabel metal2 s 77362 -960 77474 480 0 FreeSans 448 90 0 0 wbs_dat_i[18]
port 584 nsew signal input
flabel metal2 s 80858 -960 80970 480 0 FreeSans 448 90 0 0 wbs_dat_i[19]
port 585 nsew signal input
flabel metal2 s 13514 -960 13626 480 0 FreeSans 448 90 0 0 wbs_dat_i[1]
port 586 nsew signal input
flabel metal2 s 84446 -960 84558 480 0 FreeSans 448 90 0 0 wbs_dat_i[20]
port 587 nsew signal input
flabel metal2 s 87942 -960 88054 480 0 FreeSans 448 90 0 0 wbs_dat_i[21]
port 588 nsew signal input
flabel metal2 s 91530 -960 91642 480 0 FreeSans 448 90 0 0 wbs_dat_i[22]
port 589 nsew signal input
flabel metal2 s 95118 -960 95230 480 0 FreeSans 448 90 0 0 wbs_dat_i[23]
port 590 nsew signal input
flabel metal2 s 98614 -960 98726 480 0 FreeSans 448 90 0 0 wbs_dat_i[24]
port 591 nsew signal input
flabel metal2 s 102202 -960 102314 480 0 FreeSans 448 90 0 0 wbs_dat_i[25]
port 592 nsew signal input
flabel metal2 s 105698 -960 105810 480 0 FreeSans 448 90 0 0 wbs_dat_i[26]
port 593 nsew signal input
flabel metal2 s 109286 -960 109398 480 0 FreeSans 448 90 0 0 wbs_dat_i[27]
port 594 nsew signal input
flabel metal2 s 112782 -960 112894 480 0 FreeSans 448 90 0 0 wbs_dat_i[28]
port 595 nsew signal input
flabel metal2 s 116370 -960 116482 480 0 FreeSans 448 90 0 0 wbs_dat_i[29]
port 596 nsew signal input
flabel metal2 s 18206 -960 18318 480 0 FreeSans 448 90 0 0 wbs_dat_i[2]
port 597 nsew signal input
flabel metal2 s 119866 -960 119978 480 0 FreeSans 448 90 0 0 wbs_dat_i[30]
port 598 nsew signal input
flabel metal2 s 123454 -960 123566 480 0 FreeSans 448 90 0 0 wbs_dat_i[31]
port 599 nsew signal input
flabel metal2 s 22990 -960 23102 480 0 FreeSans 448 90 0 0 wbs_dat_i[3]
port 600 nsew signal input
flabel metal2 s 27682 -960 27794 480 0 FreeSans 448 90 0 0 wbs_dat_i[4]
port 601 nsew signal input
flabel metal2 s 31270 -960 31382 480 0 FreeSans 448 90 0 0 wbs_dat_i[5]
port 602 nsew signal input
flabel metal2 s 34766 -960 34878 480 0 FreeSans 448 90 0 0 wbs_dat_i[6]
port 603 nsew signal input
flabel metal2 s 38354 -960 38466 480 0 FreeSans 448 90 0 0 wbs_dat_i[7]
port 604 nsew signal input
flabel metal2 s 41850 -960 41962 480 0 FreeSans 448 90 0 0 wbs_dat_i[8]
port 605 nsew signal input
flabel metal2 s 45438 -960 45550 480 0 FreeSans 448 90 0 0 wbs_dat_i[9]
port 606 nsew signal input
flabel metal2 s 9926 -960 10038 480 0 FreeSans 448 90 0 0 wbs_dat_o[0]
port 607 nsew signal tristate
flabel metal2 s 50130 -960 50242 480 0 FreeSans 448 90 0 0 wbs_dat_o[10]
port 608 nsew signal tristate
flabel metal2 s 53718 -960 53830 480 0 FreeSans 448 90 0 0 wbs_dat_o[11]
port 609 nsew signal tristate
flabel metal2 s 57214 -960 57326 480 0 FreeSans 448 90 0 0 wbs_dat_o[12]
port 610 nsew signal tristate
flabel metal2 s 60802 -960 60914 480 0 FreeSans 448 90 0 0 wbs_dat_o[13]
port 611 nsew signal tristate
flabel metal2 s 64298 -960 64410 480 0 FreeSans 448 90 0 0 wbs_dat_o[14]
port 612 nsew signal tristate
flabel metal2 s 67886 -960 67998 480 0 FreeSans 448 90 0 0 wbs_dat_o[15]
port 613 nsew signal tristate
flabel metal2 s 71474 -960 71586 480 0 FreeSans 448 90 0 0 wbs_dat_o[16]
port 614 nsew signal tristate
flabel metal2 s 74970 -960 75082 480 0 FreeSans 448 90 0 0 wbs_dat_o[17]
port 615 nsew signal tristate
flabel metal2 s 78558 -960 78670 480 0 FreeSans 448 90 0 0 wbs_dat_o[18]
port 616 nsew signal tristate
flabel metal2 s 82054 -960 82166 480 0 FreeSans 448 90 0 0 wbs_dat_o[19]
port 617 nsew signal tristate
flabel metal2 s 14710 -960 14822 480 0 FreeSans 448 90 0 0 wbs_dat_o[1]
port 618 nsew signal tristate
flabel metal2 s 85642 -960 85754 480 0 FreeSans 448 90 0 0 wbs_dat_o[20]
port 619 nsew signal tristate
flabel metal2 s 89138 -960 89250 480 0 FreeSans 448 90 0 0 wbs_dat_o[21]
port 620 nsew signal tristate
flabel metal2 s 92726 -960 92838 480 0 FreeSans 448 90 0 0 wbs_dat_o[22]
port 621 nsew signal tristate
flabel metal2 s 96222 -960 96334 480 0 FreeSans 448 90 0 0 wbs_dat_o[23]
port 622 nsew signal tristate
flabel metal2 s 99810 -960 99922 480 0 FreeSans 448 90 0 0 wbs_dat_o[24]
port 623 nsew signal tristate
flabel metal2 s 103306 -960 103418 480 0 FreeSans 448 90 0 0 wbs_dat_o[25]
port 624 nsew signal tristate
flabel metal2 s 106894 -960 107006 480 0 FreeSans 448 90 0 0 wbs_dat_o[26]
port 625 nsew signal tristate
flabel metal2 s 110482 -960 110594 480 0 FreeSans 448 90 0 0 wbs_dat_o[27]
port 626 nsew signal tristate
flabel metal2 s 113978 -960 114090 480 0 FreeSans 448 90 0 0 wbs_dat_o[28]
port 627 nsew signal tristate
flabel metal2 s 117566 -960 117678 480 0 FreeSans 448 90 0 0 wbs_dat_o[29]
port 628 nsew signal tristate
flabel metal2 s 19402 -960 19514 480 0 FreeSans 448 90 0 0 wbs_dat_o[2]
port 629 nsew signal tristate
flabel metal2 s 121062 -960 121174 480 0 FreeSans 448 90 0 0 wbs_dat_o[30]
port 630 nsew signal tristate
flabel metal2 s 124650 -960 124762 480 0 FreeSans 448 90 0 0 wbs_dat_o[31]
port 631 nsew signal tristate
flabel metal2 s 24186 -960 24298 480 0 FreeSans 448 90 0 0 wbs_dat_o[3]
port 632 nsew signal tristate
flabel metal2 s 28878 -960 28990 480 0 FreeSans 448 90 0 0 wbs_dat_o[4]
port 633 nsew signal tristate
flabel metal2 s 32374 -960 32486 480 0 FreeSans 448 90 0 0 wbs_dat_o[5]
port 634 nsew signal tristate
flabel metal2 s 35962 -960 36074 480 0 FreeSans 448 90 0 0 wbs_dat_o[6]
port 635 nsew signal tristate
flabel metal2 s 39550 -960 39662 480 0 FreeSans 448 90 0 0 wbs_dat_o[7]
port 636 nsew signal tristate
flabel metal2 s 43046 -960 43158 480 0 FreeSans 448 90 0 0 wbs_dat_o[8]
port 637 nsew signal tristate
flabel metal2 s 46634 -960 46746 480 0 FreeSans 448 90 0 0 wbs_dat_o[9]
port 638 nsew signal tristate
flabel metal2 s 11122 -960 11234 480 0 FreeSans 448 90 0 0 wbs_sel_i[0]
port 639 nsew signal input
flabel metal2 s 15906 -960 16018 480 0 FreeSans 448 90 0 0 wbs_sel_i[1]
port 640 nsew signal input
flabel metal2 s 20598 -960 20710 480 0 FreeSans 448 90 0 0 wbs_sel_i[2]
port 641 nsew signal input
flabel metal2 s 25290 -960 25402 480 0 FreeSans 448 90 0 0 wbs_sel_i[3]
port 642 nsew signal input
flabel metal2 s 5234 -960 5346 480 0 FreeSans 448 90 0 0 wbs_stb_i
port 643 nsew signal input
flabel metal2 s 6430 -960 6542 480 0 FreeSans 448 90 0 0 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
