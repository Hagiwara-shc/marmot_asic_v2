magic
tech sky130B
magscale 1 2
timestamp 1661762021
<< metal1 >>
rect 186498 702992 186504 703044
rect 186556 703032 186562 703044
rect 188430 703032 188436 703044
rect 186556 703004 188436 703032
rect 186556 702992 186562 703004
rect 188430 702992 188436 703004
rect 188488 702992 188494 703044
rect 235166 702992 235172 703044
rect 235224 703032 235230 703044
rect 236178 703032 236184 703044
rect 235224 703004 236184 703032
rect 235224 702992 235230 703004
rect 236178 702992 236184 703004
rect 236236 702992 236242 703044
rect 522758 702992 522764 703044
rect 522816 703032 522822 703044
rect 527082 703032 527088 703044
rect 522816 703004 527088 703032
rect 522816 702992 522822 703004
rect 527082 702992 527088 703004
rect 527140 702992 527146 703044
rect 570506 702992 570512 703044
rect 570564 703032 570570 703044
rect 575842 703032 575848 703044
rect 570564 703004 575848 703032
rect 570564 702992 570570 703004
rect 575842 702992 575848 703004
rect 575900 702992 575906 703044
rect 490926 702720 490932 702772
rect 490984 702760 490990 702772
rect 494790 702760 494796 702772
rect 490984 702732 494796 702760
rect 490984 702720 490990 702732
rect 494790 702720 494796 702732
rect 494848 702720 494854 702772
rect 538674 702720 538680 702772
rect 538732 702760 538738 702772
rect 543458 702760 543464 702772
rect 538732 702732 543464 702760
rect 538732 702720 538738 702732
rect 543458 702720 543464 702732
rect 543516 702720 543522 702772
rect 24302 702448 24308 702500
rect 24360 702488 24366 702500
rect 29270 702488 29276 702500
rect 24360 702460 29276 702488
rect 24360 702448 24366 702460
rect 29270 702448 29276 702460
rect 29328 702448 29334 702500
rect 218974 702448 218980 702500
rect 219032 702488 219038 702500
rect 220262 702488 220268 702500
rect 219032 702460 220268 702488
rect 219032 702448 219038 702460
rect 220262 702448 220268 702460
rect 220320 702448 220326 702500
rect 459094 702448 459100 702500
rect 459152 702488 459158 702500
rect 462314 702488 462320 702500
rect 459152 702460 462320 702488
rect 459152 702448 459158 702460
rect 462314 702448 462320 702460
rect 462372 702448 462378 702500
rect 506842 702448 506848 702500
rect 506900 702488 506906 702500
rect 510982 702488 510988 702500
rect 506900 702460 510988 702488
rect 506900 702448 506906 702460
rect 510982 702448 510988 702460
rect 511040 702448 511046 702500
rect 554590 702448 554596 702500
rect 554648 702488 554654 702500
rect 559650 702488 559656 702500
rect 554648 702460 559656 702488
rect 554648 702448 554654 702460
rect 559650 702448 559656 702460
rect 559708 702448 559714 702500
rect 8110 700952 8116 701004
rect 8168 700992 8174 701004
rect 13078 700992 13084 701004
rect 8168 700964 13084 700992
rect 8168 700952 8174 700964
rect 13078 700952 13084 700964
rect 13136 700952 13142 701004
rect 40494 700952 40500 701004
rect 40552 700992 40558 701004
rect 44910 700992 44916 701004
rect 40552 700964 44916 700992
rect 40552 700952 40558 700964
rect 44910 700952 44916 700964
rect 44968 700952 44974 701004
rect 56778 700952 56784 701004
rect 56836 700992 56842 701004
rect 60734 700992 60740 701004
rect 56836 700964 60740 700992
rect 56836 700952 56842 700964
rect 60734 700952 60740 700964
rect 60792 700952 60798 701004
rect 72970 700952 72976 701004
rect 73028 700992 73034 701004
rect 76742 700992 76748 701004
rect 73028 700964 76748 700992
rect 73028 700952 73034 700964
rect 76742 700952 76748 700964
rect 76800 700952 76806 701004
rect 89162 700952 89168 701004
rect 89220 700992 89226 701004
rect 92566 700992 92572 701004
rect 89220 700964 92572 700992
rect 89220 700952 89226 700964
rect 92566 700952 92572 700964
rect 92624 700952 92630 701004
rect 105446 700952 105452 701004
rect 105504 700992 105510 701004
rect 108574 700992 108580 701004
rect 105504 700964 108580 700992
rect 105504 700952 105510 700964
rect 108574 700952 108580 700964
rect 108632 700952 108638 701004
rect 121638 700952 121644 701004
rect 121696 700992 121702 701004
rect 124398 700992 124404 701004
rect 121696 700964 124404 700992
rect 121696 700952 121702 700964
rect 124398 700952 124404 700964
rect 124456 700952 124462 701004
rect 137830 700952 137836 701004
rect 137888 700992 137894 701004
rect 140406 700992 140412 701004
rect 137888 700964 140412 700992
rect 137888 700952 137894 700964
rect 140406 700952 140412 700964
rect 140464 700952 140470 701004
rect 154114 700952 154120 701004
rect 154172 700992 154178 701004
rect 156230 700992 156236 701004
rect 154172 700964 156236 700992
rect 154172 700952 154178 700964
rect 156230 700952 156236 700964
rect 156288 700952 156294 701004
rect 170306 700952 170312 701004
rect 170364 700992 170370 701004
rect 172422 700992 172428 701004
rect 170364 700964 172428 700992
rect 170364 700952 170370 700964
rect 172422 700952 172428 700964
rect 172480 700952 172486 701004
rect 202782 700952 202788 701004
rect 202840 700992 202846 701004
rect 204254 700992 204260 701004
rect 202840 700964 204260 700992
rect 202840 700952 202846 700964
rect 204254 700952 204260 700964
rect 204312 700952 204318 701004
rect 348050 700952 348056 701004
rect 348108 700992 348114 701004
rect 348786 700992 348792 701004
rect 348108 700964 348792 700992
rect 348108 700952 348114 700964
rect 348786 700952 348792 700964
rect 348844 700952 348850 701004
rect 363874 700952 363880 701004
rect 363932 700992 363938 701004
rect 364978 700992 364984 701004
rect 363932 700964 364984 700992
rect 363932 700952 363938 700964
rect 364978 700952 364984 700964
rect 365036 700952 365042 701004
rect 379330 700952 379336 701004
rect 379388 700992 379394 701004
rect 381170 700992 381176 701004
rect 379388 700964 381176 700992
rect 379388 700952 379394 700964
rect 381170 700952 381176 700964
rect 381228 700952 381234 701004
rect 395706 700952 395712 701004
rect 395764 700992 395770 701004
rect 397454 700992 397460 701004
rect 395764 700964 397460 700992
rect 395764 700952 395770 700964
rect 397454 700952 397460 700964
rect 397512 700952 397518 701004
rect 411714 700952 411720 701004
rect 411772 700992 411778 701004
rect 413646 700992 413652 701004
rect 411772 700964 413652 700992
rect 411772 700952 411778 700964
rect 413646 700952 413652 700964
rect 413704 700952 413710 701004
rect 427538 700952 427544 701004
rect 427596 700992 427602 701004
rect 429838 700992 429844 701004
rect 427596 700964 429844 700992
rect 427596 700952 427602 700964
rect 429838 700952 429844 700964
rect 429896 700952 429902 701004
rect 443546 700952 443552 701004
rect 443604 700992 443610 701004
rect 446122 700992 446128 701004
rect 443604 700964 446128 700992
rect 443604 700952 443610 700964
rect 446122 700952 446128 700964
rect 446180 700952 446186 701004
rect 475378 700952 475384 701004
rect 475436 700992 475442 701004
rect 478506 700992 478512 701004
rect 475436 700964 478512 700992
rect 475436 700952 475442 700964
rect 478506 700952 478512 700964
rect 478564 700952 478570 701004
rect 74718 3992 74724 4004
rect 60706 3964 74724 3992
rect 59722 3816 59728 3868
rect 59780 3856 59786 3868
rect 60706 3856 60734 3964
rect 74718 3952 74724 3964
rect 74776 3952 74782 4004
rect 70210 3924 70216 3936
rect 59780 3828 60734 3856
rect 61856 3896 70216 3924
rect 59780 3816 59786 3828
rect 58802 3680 58808 3732
rect 58860 3720 58866 3732
rect 61856 3720 61884 3896
rect 70210 3884 70216 3896
rect 70268 3884 70274 3936
rect 78030 3924 78036 3936
rect 76392 3896 78036 3924
rect 62022 3748 62028 3800
rect 62080 3788 62086 3800
rect 67450 3788 67456 3800
rect 62080 3760 67456 3788
rect 62080 3748 62086 3760
rect 67450 3748 67456 3760
rect 67508 3748 67514 3800
rect 76392 3788 76420 3896
rect 78030 3884 78036 3896
rect 78088 3884 78094 3936
rect 83550 3856 83556 3868
rect 67560 3760 76420 3788
rect 77496 3828 83556 3856
rect 58860 3692 61884 3720
rect 58860 3680 58866 3692
rect 63218 3612 63224 3664
rect 63276 3652 63282 3664
rect 67560 3652 67588 3760
rect 69014 3680 69020 3732
rect 69072 3720 69078 3732
rect 71406 3720 71412 3732
rect 69072 3692 71412 3720
rect 69072 3680 69078 3692
rect 71406 3680 71412 3692
rect 71464 3680 71470 3732
rect 63276 3624 67588 3652
rect 63276 3612 63282 3624
rect 69106 3612 69112 3664
rect 69164 3652 69170 3664
rect 77496 3652 77524 3828
rect 83550 3816 83556 3828
rect 83608 3816 83614 3868
rect 94590 3856 94596 3868
rect 84166 3828 94596 3856
rect 80882 3748 80888 3800
rect 80940 3788 80946 3800
rect 84166 3788 84194 3828
rect 94590 3816 94596 3828
rect 94648 3816 94654 3868
rect 122282 3816 122288 3868
rect 122340 3856 122346 3868
rect 133230 3856 133236 3868
rect 122340 3828 133236 3856
rect 122340 3816 122346 3828
rect 133230 3816 133236 3828
rect 133288 3816 133294 3868
rect 80940 3760 84194 3788
rect 80940 3748 80946 3760
rect 84470 3748 84476 3800
rect 84528 3788 84534 3800
rect 97994 3788 98000 3800
rect 84528 3760 98000 3788
rect 84528 3748 84534 3760
rect 97994 3748 98000 3760
rect 98052 3748 98058 3800
rect 114002 3748 114008 3800
rect 114060 3788 114066 3800
rect 125502 3788 125508 3800
rect 114060 3760 125508 3788
rect 114060 3748 114066 3760
rect 125502 3748 125508 3760
rect 125560 3748 125566 3800
rect 81342 3720 81348 3732
rect 69164 3624 77524 3652
rect 77588 3692 81348 3720
rect 69164 3612 69170 3624
rect 66714 3544 66720 3596
rect 66772 3584 66778 3596
rect 77588 3584 77616 3692
rect 81342 3680 81348 3692
rect 81400 3680 81406 3732
rect 85666 3680 85672 3732
rect 85724 3720 85730 3732
rect 85724 3692 87000 3720
rect 85724 3680 85730 3692
rect 86862 3652 86868 3664
rect 66772 3556 77616 3584
rect 77680 3624 86868 3652
rect 66772 3544 66778 3556
rect 56042 3476 56048 3528
rect 56100 3516 56106 3528
rect 69014 3516 69020 3528
rect 56100 3488 69020 3516
rect 56100 3476 56106 3488
rect 69014 3476 69020 3488
rect 69072 3476 69078 3528
rect 70118 3476 70124 3528
rect 70176 3516 70182 3528
rect 70176 3488 70394 3516
rect 70176 3476 70182 3488
rect 54938 3408 54944 3460
rect 54996 3448 55002 3460
rect 70210 3448 70216 3460
rect 54996 3420 70216 3448
rect 54996 3408 55002 3420
rect 70210 3408 70216 3420
rect 70268 3408 70274 3460
rect 70366 3448 70394 3488
rect 72970 3476 72976 3528
rect 73028 3516 73034 3528
rect 77680 3516 77708 3624
rect 86862 3612 86868 3624
rect 86920 3612 86926 3664
rect 86972 3652 87000 3692
rect 87782 3680 87788 3732
rect 87840 3720 87846 3732
rect 101214 3720 101220 3732
rect 87840 3692 101220 3720
rect 87840 3680 87846 3692
rect 101214 3680 101220 3692
rect 101272 3680 101278 3732
rect 116394 3680 116400 3732
rect 116452 3720 116458 3732
rect 127710 3720 127716 3732
rect 116452 3692 127716 3720
rect 116452 3680 116458 3692
rect 127710 3680 127716 3692
rect 127768 3680 127774 3732
rect 99006 3652 99012 3664
rect 86972 3624 99012 3652
rect 99006 3612 99012 3624
rect 99064 3612 99070 3664
rect 109402 3612 109408 3664
rect 109460 3652 109466 3664
rect 121178 3652 121184 3664
rect 109460 3624 121184 3652
rect 109460 3612 109466 3624
rect 121178 3612 121184 3624
rect 121236 3612 121242 3664
rect 125042 3612 125048 3664
rect 125100 3652 125106 3664
rect 135438 3652 135444 3664
rect 125100 3624 135444 3652
rect 125100 3612 125106 3624
rect 135438 3612 135444 3624
rect 135496 3612 135502 3664
rect 143626 3612 143632 3664
rect 143684 3652 143690 3664
rect 153102 3652 153108 3664
rect 143684 3624 153108 3652
rect 143684 3612 143690 3624
rect 153102 3612 153108 3624
rect 153160 3612 153166 3664
rect 82906 3584 82912 3596
rect 73028 3488 77708 3516
rect 78508 3556 82912 3584
rect 73028 3476 73034 3488
rect 78508 3448 78536 3556
rect 82906 3544 82912 3556
rect 82964 3544 82970 3596
rect 83274 3544 83280 3596
rect 83332 3584 83338 3596
rect 96798 3584 96804 3596
rect 83332 3556 96804 3584
rect 83332 3544 83338 3556
rect 96798 3544 96804 3556
rect 96856 3544 96862 3596
rect 102226 3544 102232 3596
rect 102284 3584 102290 3596
rect 114462 3584 114468 3596
rect 102284 3556 114468 3584
rect 102284 3544 102290 3556
rect 114462 3544 114468 3556
rect 114520 3544 114526 3596
rect 121086 3544 121092 3596
rect 121144 3584 121150 3596
rect 132126 3584 132132 3596
rect 121144 3556 132132 3584
rect 121144 3544 121150 3556
rect 132126 3544 132132 3556
rect 132184 3544 132190 3596
rect 136450 3544 136456 3596
rect 136508 3584 136514 3596
rect 146478 3584 146484 3596
rect 136508 3556 146484 3584
rect 136508 3544 136514 3556
rect 146478 3544 146484 3556
rect 146536 3544 146542 3596
rect 149514 3544 149520 3596
rect 149572 3584 149578 3596
rect 158622 3584 158628 3596
rect 149572 3556 158628 3584
rect 149572 3544 149578 3556
rect 158622 3544 158628 3556
rect 158680 3544 158686 3596
rect 78582 3476 78588 3528
rect 78640 3516 78646 3528
rect 92382 3516 92388 3528
rect 78640 3488 92388 3516
rect 78640 3476 78646 3488
rect 92382 3476 92388 3488
rect 92440 3476 92446 3528
rect 103606 3516 103612 3528
rect 92492 3488 103612 3516
rect 85758 3448 85764 3460
rect 70366 3420 78536 3448
rect 79428 3420 85764 3448
rect 51350 3340 51356 3392
rect 51408 3380 51414 3392
rect 66990 3380 66996 3392
rect 51408 3352 66996 3380
rect 51408 3340 51414 3352
rect 66990 3340 66996 3352
rect 67048 3340 67054 3392
rect 67450 3340 67456 3392
rect 67508 3380 67514 3392
rect 76926 3380 76932 3392
rect 67508 3352 76932 3380
rect 67508 3340 67514 3352
rect 76926 3340 76932 3352
rect 76984 3340 76990 3392
rect 65518 3272 65524 3324
rect 65576 3312 65582 3324
rect 65576 3284 70394 3312
rect 65576 3272 65582 3284
rect 50154 3204 50160 3256
rect 50212 3244 50218 3256
rect 65886 3244 65892 3256
rect 50212 3216 65892 3244
rect 50212 3204 50218 3216
rect 65886 3204 65892 3216
rect 65944 3204 65950 3256
rect 70366 3244 70394 3284
rect 71498 3272 71504 3324
rect 71556 3312 71562 3324
rect 79428 3312 79456 3420
rect 85758 3408 85764 3420
rect 85816 3408 85822 3460
rect 90358 3408 90364 3460
rect 90416 3448 90422 3460
rect 92492 3448 92520 3488
rect 103606 3476 103612 3488
rect 103664 3476 103670 3528
rect 110506 3476 110512 3528
rect 110564 3516 110570 3528
rect 122374 3516 122380 3528
rect 110564 3488 122380 3516
rect 110564 3476 110570 3488
rect 122374 3476 122380 3488
rect 122432 3476 122438 3528
rect 127066 3476 127072 3528
rect 127124 3516 127130 3528
rect 137646 3516 137652 3528
rect 127124 3488 137652 3516
rect 127124 3476 127130 3488
rect 137646 3476 137652 3488
rect 137704 3476 137710 3528
rect 139210 3476 139216 3528
rect 139268 3516 139274 3528
rect 148686 3516 148692 3528
rect 139268 3488 148692 3516
rect 139268 3476 139274 3488
rect 148686 3476 148692 3488
rect 148744 3476 148750 3528
rect 153010 3476 153016 3528
rect 153068 3516 153074 3528
rect 160186 3516 160192 3528
rect 153068 3488 160192 3516
rect 153068 3476 153074 3488
rect 160186 3476 160192 3488
rect 160244 3476 160250 3528
rect 102318 3448 102324 3460
rect 90416 3420 92520 3448
rect 93826 3420 102324 3448
rect 90416 3408 90422 3420
rect 79686 3340 79692 3392
rect 79744 3380 79750 3392
rect 82998 3380 83004 3392
rect 79744 3352 83004 3380
rect 79744 3340 79750 3352
rect 82998 3340 83004 3352
rect 83056 3340 83062 3392
rect 89530 3340 89536 3392
rect 89588 3380 89594 3392
rect 93826 3380 93854 3420
rect 102318 3408 102324 3420
rect 102376 3408 102382 3460
rect 105722 3408 105728 3460
rect 105780 3448 105786 3460
rect 117774 3448 117780 3460
rect 105780 3420 117780 3448
rect 105780 3408 105786 3420
rect 117774 3408 117780 3420
rect 117832 3408 117838 3460
rect 131758 3408 131764 3460
rect 131816 3448 131822 3460
rect 142246 3448 142252 3460
rect 131816 3420 142252 3448
rect 131816 3408 131822 3420
rect 142246 3408 142252 3420
rect 142304 3408 142310 3460
rect 142522 3408 142528 3460
rect 142580 3448 142586 3460
rect 151722 3448 151728 3460
rect 142580 3420 151728 3448
rect 142580 3408 142586 3420
rect 151722 3408 151728 3420
rect 151780 3408 151786 3460
rect 155770 3408 155776 3460
rect 155828 3448 155834 3460
rect 155828 3420 157380 3448
rect 155828 3408 155834 3420
rect 89588 3352 93854 3380
rect 89588 3340 89594 3352
rect 96246 3340 96252 3392
rect 96304 3380 96310 3392
rect 109034 3380 109040 3392
rect 96304 3352 109040 3380
rect 96304 3340 96310 3352
rect 109034 3340 109040 3352
rect 109092 3340 109098 3392
rect 112806 3340 112812 3392
rect 112864 3380 112870 3392
rect 124122 3380 124128 3392
rect 112864 3352 124128 3380
rect 112864 3340 112870 3352
rect 124122 3340 124128 3352
rect 124180 3340 124186 3392
rect 125962 3340 125968 3392
rect 126020 3380 126026 3392
rect 136634 3380 136640 3392
rect 126020 3352 136640 3380
rect 126020 3340 126026 3352
rect 136634 3340 136640 3352
rect 136692 3340 136698 3392
rect 149790 3380 149796 3392
rect 140056 3352 149796 3380
rect 71556 3284 79456 3312
rect 71556 3272 71562 3284
rect 82906 3272 82912 3324
rect 82964 3312 82970 3324
rect 84654 3312 84660 3324
rect 82964 3284 84660 3312
rect 82964 3272 82970 3284
rect 84654 3272 84660 3284
rect 84712 3272 84718 3324
rect 86862 3272 86868 3324
rect 86920 3312 86926 3324
rect 100110 3312 100116 3324
rect 86920 3284 100116 3312
rect 86920 3272 86926 3284
rect 100110 3272 100116 3284
rect 100168 3272 100174 3324
rect 103330 3272 103336 3324
rect 103388 3312 103394 3324
rect 115566 3312 115572 3324
rect 103388 3284 115572 3312
rect 103388 3272 103394 3284
rect 115566 3272 115572 3284
rect 115624 3272 115630 3324
rect 117590 3272 117596 3324
rect 117648 3312 117654 3324
rect 128814 3312 128820 3324
rect 117648 3284 128820 3312
rect 117648 3272 117654 3284
rect 128814 3272 128820 3284
rect 128872 3272 128878 3324
rect 129366 3272 129372 3324
rect 129424 3312 129430 3324
rect 139854 3312 139860 3324
rect 129424 3284 139860 3312
rect 129424 3272 129430 3284
rect 139854 3272 139860 3284
rect 139912 3272 139918 3324
rect 140056 3256 140084 3352
rect 149790 3340 149796 3352
rect 149848 3340 149854 3392
rect 148318 3272 148324 3324
rect 148376 3312 148382 3324
rect 157242 3312 157248 3324
rect 148376 3284 157248 3312
rect 148376 3272 148382 3284
rect 157242 3272 157248 3284
rect 157300 3272 157306 3324
rect 79962 3244 79968 3256
rect 70366 3216 79968 3244
rect 79962 3204 79968 3216
rect 80020 3204 80026 3256
rect 93946 3204 93952 3256
rect 94004 3244 94010 3256
rect 106734 3244 106740 3256
rect 94004 3216 106740 3244
rect 94004 3204 94010 3216
rect 106734 3204 106740 3216
rect 106792 3204 106798 3256
rect 107194 3204 107200 3256
rect 107252 3244 107258 3256
rect 118602 3244 118608 3256
rect 107252 3216 118608 3244
rect 107252 3204 107258 3216
rect 118602 3204 118608 3216
rect 118660 3204 118666 3256
rect 119890 3204 119896 3256
rect 119948 3244 119954 3256
rect 131022 3244 131028 3256
rect 119948 3216 131028 3244
rect 119948 3204 119954 3216
rect 131022 3204 131028 3216
rect 131080 3204 131086 3256
rect 140038 3204 140044 3256
rect 140096 3204 140102 3256
rect 154022 3204 154028 3256
rect 154080 3244 154086 3256
rect 154080 3216 156552 3244
rect 154080 3204 154086 3216
rect 40954 3136 40960 3188
rect 41012 3176 41018 3188
rect 57054 3176 57060 3188
rect 41012 3148 57060 3176
rect 41012 3136 41018 3148
rect 57054 3136 57060 3148
rect 57112 3136 57118 3188
rect 57514 3136 57520 3188
rect 57572 3176 57578 3188
rect 72510 3176 72516 3188
rect 57572 3148 72516 3176
rect 57572 3136 57578 3148
rect 72510 3136 72516 3148
rect 72568 3136 72574 3188
rect 73798 3136 73804 3188
rect 73856 3176 73862 3188
rect 87966 3176 87972 3188
rect 73856 3148 87972 3176
rect 73856 3136 73862 3148
rect 87966 3136 87972 3148
rect 88024 3136 88030 3188
rect 101030 3136 101036 3188
rect 101088 3176 101094 3188
rect 113082 3176 113088 3188
rect 101088 3148 113088 3176
rect 101088 3136 101094 3148
rect 113082 3136 113088 3148
rect 113140 3136 113146 3188
rect 134334 3176 134340 3188
rect 123496 3148 134340 3176
rect 52546 3068 52552 3120
rect 52604 3108 52610 3120
rect 68094 3108 68100 3120
rect 52604 3080 68100 3108
rect 52604 3068 52610 3080
rect 68094 3068 68100 3080
rect 68152 3068 68158 3120
rect 76282 3068 76288 3120
rect 76340 3108 76346 3120
rect 76340 3080 79272 3108
rect 76340 3068 76346 3080
rect 44266 3000 44272 3052
rect 44324 3040 44330 3052
rect 60366 3040 60372 3052
rect 44324 3012 60372 3040
rect 44324 3000 44330 3012
rect 60366 3000 60372 3012
rect 60424 3000 60430 3052
rect 64322 3000 64328 3052
rect 64380 3040 64386 3052
rect 79134 3040 79140 3052
rect 64380 3012 79140 3040
rect 64380 3000 64386 3012
rect 79134 3000 79140 3012
rect 79192 3000 79198 3052
rect 79244 3040 79272 3080
rect 79594 3068 79600 3120
rect 79652 3108 79658 3120
rect 89070 3108 89076 3120
rect 79652 3080 89076 3108
rect 79652 3068 79658 3080
rect 89070 3068 89076 3080
rect 89128 3068 89134 3120
rect 98730 3068 98736 3120
rect 98788 3108 98794 3120
rect 111150 3108 111156 3120
rect 98788 3080 111156 3108
rect 98788 3068 98794 3080
rect 111150 3068 111156 3080
rect 111208 3068 111214 3120
rect 111610 3068 111616 3120
rect 111668 3108 111674 3120
rect 123294 3108 123300 3120
rect 111668 3080 123300 3108
rect 111668 3068 111674 3080
rect 123294 3068 123300 3080
rect 123352 3068 123358 3120
rect 79244 3012 82860 3040
rect 33594 2932 33600 2984
rect 33652 2972 33658 2984
rect 50430 2972 50436 2984
rect 33652 2944 50436 2972
rect 33652 2932 33658 2944
rect 50430 2932 50436 2944
rect 50488 2932 50494 2984
rect 64874 2972 64880 2984
rect 50632 2944 64880 2972
rect 26602 2864 26608 2916
rect 26660 2904 26666 2916
rect 43806 2904 43812 2916
rect 26660 2876 43812 2904
rect 26660 2864 26666 2876
rect 43806 2864 43812 2876
rect 43864 2864 43870 2916
rect 48958 2864 48964 2916
rect 49016 2904 49022 2916
rect 50632 2904 50660 2944
rect 64874 2932 64880 2944
rect 64932 2932 64938 2984
rect 67910 2932 67916 2984
rect 67968 2972 67974 2984
rect 82722 2972 82728 2984
rect 67968 2944 82728 2972
rect 67968 2932 67974 2944
rect 82722 2932 82728 2944
rect 82780 2932 82786 2984
rect 82832 2972 82860 3012
rect 82998 3000 83004 3052
rect 83056 3040 83062 3052
rect 93486 3040 93492 3052
rect 83056 3012 93492 3040
rect 83056 3000 83062 3012
rect 93486 3000 93492 3012
rect 93544 3000 93550 3052
rect 95142 3000 95148 3052
rect 95200 3040 95206 3052
rect 107838 3040 107844 3052
rect 95200 3012 107844 3040
rect 95200 3000 95206 3012
rect 107838 3000 107844 3012
rect 107896 3000 107902 3052
rect 108482 3000 108488 3052
rect 108540 3040 108546 3052
rect 119982 3040 119988 3052
rect 108540 3012 119988 3040
rect 108540 3000 108546 3012
rect 119982 3000 119988 3012
rect 120040 3000 120046 3052
rect 123496 2984 123524 3148
rect 134334 3136 134340 3148
rect 134392 3136 134398 3188
rect 137646 3136 137652 3188
rect 137704 3176 137710 3188
rect 147766 3176 147772 3188
rect 137704 3148 147772 3176
rect 137704 3136 137710 3148
rect 147766 3136 147772 3148
rect 147824 3136 147830 3188
rect 156414 3176 156420 3188
rect 151556 3148 156420 3176
rect 134150 3068 134156 3120
rect 134208 3108 134214 3120
rect 144270 3108 144276 3120
rect 134208 3080 144276 3108
rect 134208 3068 134214 3080
rect 144270 3068 144276 3080
rect 144328 3068 144334 3120
rect 147122 3068 147128 3120
rect 147180 3108 147186 3120
rect 151556 3108 151584 3148
rect 156414 3136 156420 3148
rect 156472 3136 156478 3188
rect 155310 3108 155316 3120
rect 147180 3080 151584 3108
rect 151648 3080 155316 3108
rect 147180 3068 147186 3080
rect 128170 3000 128176 3052
rect 128228 3040 128234 3052
rect 138750 3040 138756 3052
rect 128228 3012 138756 3040
rect 128228 3000 128234 3012
rect 138750 3000 138756 3012
rect 138808 3000 138814 3052
rect 143166 3040 143172 3052
rect 141068 3012 143172 3040
rect 90450 2972 90456 2984
rect 82832 2944 90456 2972
rect 90450 2932 90456 2944
rect 90508 2932 90514 2984
rect 91554 2932 91560 2984
rect 91612 2972 91618 2984
rect 104526 2972 104532 2984
rect 91612 2944 104532 2972
rect 91612 2932 91618 2944
rect 104526 2932 104532 2944
rect 104584 2932 104590 2984
rect 104618 2932 104624 2984
rect 104676 2972 104682 2984
rect 116946 2972 116952 2984
rect 104676 2944 116952 2972
rect 104676 2932 104682 2944
rect 116946 2932 116952 2944
rect 117004 2932 117010 2984
rect 123478 2932 123484 2984
rect 123536 2932 123542 2984
rect 130562 2932 130568 2984
rect 130620 2972 130626 2984
rect 140958 2972 140964 2984
rect 130620 2944 140964 2972
rect 130620 2932 130626 2944
rect 140958 2932 140964 2944
rect 141016 2932 141022 2984
rect 63678 2904 63684 2916
rect 49016 2876 50660 2904
rect 55186 2876 63684 2904
rect 49016 2864 49022 2876
rect 27706 2796 27712 2848
rect 27764 2836 27770 2848
rect 45186 2836 45192 2848
rect 27764 2808 45192 2836
rect 27764 2796 27770 2808
rect 45186 2796 45192 2808
rect 45244 2796 45250 2848
rect 47854 2796 47860 2848
rect 47912 2836 47918 2848
rect 55186 2836 55214 2876
rect 63678 2864 63684 2876
rect 63736 2864 63742 2916
rect 75362 2864 75368 2916
rect 75420 2904 75426 2916
rect 79594 2904 79600 2916
rect 75420 2876 79600 2904
rect 75420 2864 75426 2876
rect 79594 2864 79600 2876
rect 79652 2864 79658 2916
rect 82078 2864 82084 2916
rect 82136 2904 82142 2916
rect 95970 2904 95976 2916
rect 82136 2876 95976 2904
rect 82136 2864 82142 2876
rect 95970 2864 95976 2876
rect 96028 2864 96034 2916
rect 97442 2864 97448 2916
rect 97500 2904 97506 2916
rect 110046 2904 110052 2916
rect 97500 2876 110052 2904
rect 97500 2864 97506 2876
rect 110046 2864 110052 2876
rect 110104 2864 110110 2916
rect 115198 2864 115204 2916
rect 115256 2904 115262 2916
rect 126882 2904 126888 2916
rect 115256 2876 126888 2904
rect 115256 2864 115262 2876
rect 126882 2864 126888 2876
rect 126940 2864 126946 2916
rect 132954 2864 132960 2916
rect 133012 2904 133018 2916
rect 141068 2904 141096 3012
rect 143166 3000 143172 3012
rect 143224 3000 143230 3052
rect 145926 3000 145932 3052
rect 145984 3040 145990 3052
rect 151648 3040 151676 3080
rect 155310 3068 155316 3080
rect 155368 3068 155374 3120
rect 156524 3108 156552 3216
rect 157352 3176 157380 3420
rect 166074 3408 166080 3460
rect 166132 3448 166138 3460
rect 166132 3420 171134 3448
rect 166132 3408 166138 3420
rect 166350 3380 166356 3392
rect 158732 3352 166356 3380
rect 158162 3272 158168 3324
rect 158220 3312 158226 3324
rect 158732 3312 158760 3352
rect 166350 3340 166356 3352
rect 166408 3340 166414 3392
rect 171106 3380 171134 3420
rect 174078 3380 174084 3392
rect 171106 3352 174084 3380
rect 174078 3340 174084 3352
rect 174136 3340 174142 3392
rect 158220 3284 158760 3312
rect 158220 3272 158226 3284
rect 161290 3272 161296 3324
rect 161348 3312 161354 3324
rect 169662 3312 169668 3324
rect 161348 3284 169668 3312
rect 161348 3272 161354 3284
rect 169662 3272 169668 3284
rect 169720 3272 169726 3324
rect 181806 3312 181812 3324
rect 174280 3284 181812 3312
rect 174280 3256 174308 3284
rect 181806 3272 181812 3284
rect 181864 3272 181870 3324
rect 564342 3272 564348 3324
rect 564400 3312 564406 3324
rect 583386 3312 583392 3324
rect 564400 3284 583392 3312
rect 564400 3272 564406 3284
rect 583386 3272 583392 3284
rect 583444 3272 583450 3324
rect 160186 3204 160192 3256
rect 160244 3244 160250 3256
rect 161934 3244 161940 3256
rect 160244 3216 161940 3244
rect 160244 3204 160250 3216
rect 161934 3204 161940 3216
rect 161992 3204 161998 3256
rect 163682 3204 163688 3256
rect 163740 3244 163746 3256
rect 171870 3244 171876 3256
rect 163740 3216 171876 3244
rect 163740 3204 163746 3216
rect 171870 3204 171876 3216
rect 171928 3204 171934 3256
rect 174262 3204 174268 3256
rect 174320 3204 174326 3256
rect 180886 3244 180892 3256
rect 178604 3216 180892 3244
rect 164142 3176 164148 3188
rect 157352 3148 164148 3176
rect 164142 3136 164148 3148
rect 164200 3136 164206 3188
rect 170766 3136 170772 3188
rect 170824 3176 170830 3188
rect 178494 3176 178500 3188
rect 170824 3148 178500 3176
rect 170824 3136 170830 3148
rect 178494 3136 178500 3148
rect 178552 3136 178558 3188
rect 162762 3108 162768 3120
rect 156524 3080 162768 3108
rect 162762 3068 162768 3080
rect 162820 3068 162826 3120
rect 164878 3068 164884 3120
rect 164936 3108 164942 3120
rect 172974 3108 172980 3120
rect 164936 3080 172980 3108
rect 164936 3068 164942 3080
rect 172974 3068 172980 3080
rect 173032 3068 173038 3120
rect 173434 3068 173440 3120
rect 173492 3108 173498 3120
rect 178604 3108 178632 3216
rect 180886 3204 180892 3216
rect 180944 3204 180950 3256
rect 184934 3204 184940 3256
rect 184992 3244 184998 3256
rect 184992 3216 190454 3244
rect 184992 3204 184998 3216
rect 181438 3136 181444 3188
rect 181496 3176 181502 3188
rect 188430 3176 188436 3188
rect 181496 3148 188436 3176
rect 181496 3136 181502 3148
rect 188430 3136 188436 3148
rect 188488 3136 188494 3188
rect 190426 3176 190454 3216
rect 200298 3204 200304 3256
rect 200356 3244 200362 3256
rect 206094 3244 206100 3256
rect 200356 3216 206100 3244
rect 200356 3204 200362 3216
rect 206094 3204 206100 3216
rect 206152 3204 206158 3256
rect 556706 3204 556712 3256
rect 556764 3244 556770 3256
rect 575106 3244 575112 3256
rect 556764 3216 575112 3244
rect 556764 3204 556770 3216
rect 575106 3204 575112 3216
rect 575164 3204 575170 3256
rect 191742 3176 191748 3188
rect 190426 3148 191748 3176
rect 191742 3136 191748 3148
rect 191800 3136 191806 3188
rect 195606 3136 195612 3188
rect 195664 3176 195670 3188
rect 201678 3176 201684 3188
rect 195664 3148 201684 3176
rect 195664 3136 195670 3148
rect 201678 3136 201684 3148
rect 201736 3136 201742 3188
rect 220262 3136 220268 3188
rect 220320 3176 220326 3188
rect 224862 3176 224868 3188
rect 220320 3148 224868 3176
rect 220320 3136 220326 3148
rect 224862 3136 224868 3148
rect 224920 3136 224926 3188
rect 561122 3136 561128 3188
rect 561180 3176 561186 3188
rect 579798 3176 579804 3188
rect 561180 3148 579804 3176
rect 561180 3136 561186 3148
rect 579798 3136 579804 3148
rect 579856 3136 579862 3188
rect 173492 3080 178632 3108
rect 173492 3068 173498 3080
rect 179046 3068 179052 3120
rect 179104 3108 179110 3120
rect 186314 3108 186320 3120
rect 179104 3080 186320 3108
rect 179104 3068 179110 3080
rect 186314 3068 186320 3080
rect 186372 3068 186378 3120
rect 190546 3068 190552 3120
rect 190604 3108 190610 3120
rect 197262 3108 197268 3120
rect 190604 3080 197268 3108
rect 190604 3068 190610 3080
rect 197262 3068 197268 3080
rect 197320 3068 197326 3120
rect 202690 3068 202696 3120
rect 202748 3108 202754 3120
rect 208302 3108 208308 3120
rect 202748 3080 208308 3108
rect 202748 3068 202754 3080
rect 208302 3068 208308 3080
rect 208360 3068 208366 3120
rect 209866 3068 209872 3120
rect 209924 3108 209930 3120
rect 214926 3108 214932 3120
rect 209924 3080 214932 3108
rect 209924 3068 209930 3080
rect 214926 3068 214932 3080
rect 214984 3068 214990 3120
rect 215662 3068 215668 3120
rect 215720 3108 215726 3120
rect 220446 3108 220452 3120
rect 215720 3080 220452 3108
rect 215720 3068 215726 3080
rect 220446 3068 220452 3080
rect 220504 3068 220510 3120
rect 221550 3068 221556 3120
rect 221608 3108 221614 3120
rect 225966 3108 225972 3120
rect 221608 3080 225972 3108
rect 221608 3068 221614 3080
rect 225966 3068 225972 3080
rect 226024 3068 226030 3120
rect 228726 3068 228732 3120
rect 228784 3108 228790 3120
rect 232590 3108 232596 3120
rect 228784 3080 232596 3108
rect 228784 3068 228790 3080
rect 232590 3068 232596 3080
rect 232648 3068 232654 3120
rect 239306 3068 239312 3120
rect 239364 3108 239370 3120
rect 242526 3108 242532 3120
rect 239364 3080 242532 3108
rect 239364 3068 239370 3080
rect 242526 3068 242532 3080
rect 242584 3068 242590 3120
rect 543458 3068 543464 3120
rect 543516 3108 543522 3120
rect 560478 3108 560484 3120
rect 543516 3080 560484 3108
rect 543516 3068 543522 3080
rect 560478 3068 560484 3080
rect 560536 3068 560542 3120
rect 562226 3068 562232 3120
rect 562284 3108 562290 3120
rect 580994 3108 581000 3120
rect 562284 3080 581000 3108
rect 562284 3068 562290 3080
rect 580994 3068 581000 3080
rect 581052 3068 581058 3120
rect 145984 3012 151676 3040
rect 145984 3000 145990 3012
rect 151814 3000 151820 3052
rect 151872 3040 151878 3052
rect 160830 3040 160836 3052
rect 151872 3012 160836 3040
rect 151872 3000 151878 3012
rect 160830 3000 160836 3012
rect 160888 3000 160894 3052
rect 162486 3000 162492 3052
rect 162544 3040 162550 3052
rect 170858 3040 170864 3052
rect 162544 3012 170864 3040
rect 162544 3000 162550 3012
rect 170858 3000 170864 3012
rect 170916 3000 170922 3052
rect 171962 3000 171968 3052
rect 172020 3040 172026 3052
rect 179598 3040 179604 3052
rect 172020 3012 179604 3040
rect 172020 3000 172026 3012
rect 179598 3000 179604 3012
rect 179656 3000 179662 3052
rect 182542 3000 182548 3052
rect 182600 3040 182606 3052
rect 189534 3040 189540 3052
rect 182600 3012 189540 3040
rect 182600 3000 182606 3012
rect 189534 3000 189540 3012
rect 189592 3000 189598 3052
rect 189718 3000 189724 3052
rect 189776 3040 189782 3052
rect 196158 3040 196164 3052
rect 189776 3012 196164 3040
rect 189776 3000 189782 3012
rect 196158 3000 196164 3012
rect 196216 3000 196222 3052
rect 200574 3040 200580 3052
rect 196360 3012 200580 3040
rect 141234 2932 141240 2984
rect 141292 2972 141298 2984
rect 150894 2972 150900 2984
rect 141292 2944 150900 2972
rect 141292 2932 141298 2944
rect 150894 2932 150900 2944
rect 150952 2932 150958 2984
rect 156598 2932 156604 2984
rect 156656 2972 156662 2984
rect 165522 2972 165528 2984
rect 156656 2944 165528 2972
rect 156656 2932 156662 2944
rect 165522 2932 165528 2944
rect 165580 2932 165586 2984
rect 167178 2932 167184 2984
rect 167236 2972 167242 2984
rect 175458 2972 175464 2984
rect 167236 2944 175464 2972
rect 167236 2932 167242 2944
rect 175458 2932 175464 2944
rect 175516 2932 175522 2984
rect 175826 2932 175832 2984
rect 175884 2972 175890 2984
rect 175884 2944 177804 2972
rect 175884 2932 175890 2944
rect 133012 2876 141096 2904
rect 133012 2864 133018 2876
rect 144730 2864 144736 2916
rect 144788 2904 144794 2916
rect 144788 2876 147674 2904
rect 144788 2864 144794 2876
rect 47912 2808 55214 2836
rect 47912 2796 47918 2808
rect 60826 2796 60832 2848
rect 60884 2836 60890 2848
rect 75822 2836 75828 2848
rect 60884 2808 75828 2836
rect 60884 2796 60890 2808
rect 75822 2796 75828 2808
rect 75880 2796 75886 2848
rect 77386 2796 77392 2848
rect 77444 2836 77450 2848
rect 91278 2836 91284 2848
rect 77444 2808 91284 2836
rect 77444 2796 77450 2808
rect 91278 2796 91284 2808
rect 91336 2796 91342 2848
rect 92750 2796 92756 2848
rect 92808 2836 92814 2848
rect 98638 2836 98644 2848
rect 92808 2808 98644 2836
rect 92808 2796 92814 2808
rect 98638 2796 98644 2808
rect 98696 2796 98702 2848
rect 99834 2796 99840 2848
rect 99892 2836 99898 2848
rect 112530 2836 112536 2848
rect 99892 2808 112536 2836
rect 99892 2796 99898 2808
rect 112530 2796 112536 2808
rect 112588 2796 112594 2848
rect 118786 2796 118792 2848
rect 118844 2836 118850 2848
rect 130194 2836 130200 2848
rect 118844 2808 130200 2836
rect 118844 2796 118850 2808
rect 130194 2796 130200 2808
rect 130252 2796 130258 2848
rect 135254 2796 135260 2848
rect 135312 2836 135318 2848
rect 145374 2836 145380 2848
rect 135312 2808 145380 2836
rect 135312 2796 135318 2808
rect 145374 2796 145380 2808
rect 145432 2796 145438 2848
rect 147646 2836 147674 2876
rect 150618 2864 150624 2916
rect 150676 2904 150682 2916
rect 160002 2904 160008 2916
rect 150676 2876 160008 2904
rect 150676 2864 150682 2876
rect 160002 2864 160008 2876
rect 160060 2864 160066 2916
rect 160094 2864 160100 2916
rect 160152 2904 160158 2916
rect 168834 2904 168840 2916
rect 160152 2876 168840 2904
rect 160152 2864 160158 2876
rect 168834 2864 168840 2876
rect 168892 2864 168898 2916
rect 169570 2864 169576 2916
rect 169628 2904 169634 2916
rect 177666 2904 177672 2916
rect 169628 2876 177672 2904
rect 169628 2864 169634 2876
rect 177666 2864 177672 2876
rect 177724 2864 177730 2916
rect 177776 2904 177804 2944
rect 177850 2932 177856 2984
rect 177908 2972 177914 2984
rect 185394 2972 185400 2984
rect 177908 2944 185400 2972
rect 177908 2932 177914 2944
rect 185394 2932 185400 2944
rect 185452 2932 185458 2984
rect 194410 2932 194416 2984
rect 194468 2972 194474 2984
rect 196360 2972 196388 3012
rect 200574 3000 200580 3012
rect 200632 3000 200638 3052
rect 203886 3000 203892 3052
rect 203944 3040 203950 3052
rect 209406 3040 209412 3052
rect 203944 3012 209412 3040
rect 203944 3000 203950 3012
rect 209406 3000 209412 3012
rect 209464 3000 209470 3052
rect 212166 3000 212172 3052
rect 212224 3040 212230 3052
rect 217134 3040 217140 3052
rect 212224 3012 217140 3040
rect 212224 3000 212230 3012
rect 217134 3000 217140 3012
rect 217192 3000 217198 3052
rect 219250 3000 219256 3052
rect 219308 3040 219314 3052
rect 223482 3040 223488 3052
rect 219308 3012 223488 3040
rect 219308 3000 219314 3012
rect 223482 3000 223488 3012
rect 223540 3000 223546 3052
rect 228174 3040 228180 3052
rect 223960 3012 228180 3040
rect 223960 2984 223988 3012
rect 228174 3000 228180 3012
rect 228232 3000 228238 3052
rect 229830 3000 229836 3052
rect 229888 3040 229894 3052
rect 233694 3040 233700 3052
rect 229888 3012 233700 3040
rect 229888 3000 229894 3012
rect 233694 3000 233700 3012
rect 233752 3000 233758 3052
rect 234614 3000 234620 3052
rect 234672 3040 234678 3052
rect 238110 3040 238116 3052
rect 234672 3012 238116 3040
rect 234672 3000 234678 3012
rect 238110 3000 238116 3012
rect 238168 3000 238174 3052
rect 240502 3000 240508 3052
rect 240560 3040 240566 3052
rect 243630 3040 243636 3052
rect 240560 3012 243636 3040
rect 240560 3000 240566 3012
rect 243630 3000 243636 3012
rect 243688 3000 243694 3052
rect 245194 3000 245200 3052
rect 245252 3040 245258 3052
rect 248046 3040 248052 3052
rect 245252 3012 248052 3040
rect 245252 3000 245258 3012
rect 248046 3000 248052 3012
rect 248104 3000 248110 3052
rect 248782 3000 248788 3052
rect 248840 3040 248846 3052
rect 251358 3040 251364 3052
rect 248840 3012 251364 3040
rect 248840 3000 248846 3012
rect 251358 3000 251364 3012
rect 251416 3000 251422 3052
rect 333698 3000 333704 3052
rect 333756 3040 333762 3052
rect 336274 3040 336280 3052
rect 333756 3012 336280 3040
rect 333756 3000 333762 3012
rect 336274 3000 336280 3012
rect 336332 3000 336338 3052
rect 530026 3000 530032 3052
rect 530084 3040 530090 3052
rect 546678 3040 546684 3052
rect 530084 3012 546684 3040
rect 530084 3000 530090 3012
rect 546678 3000 546684 3012
rect 546736 3000 546742 3052
rect 553302 3000 553308 3052
rect 553360 3040 553366 3052
rect 571518 3040 571524 3052
rect 553360 3012 571524 3040
rect 553360 3000 553366 3012
rect 571518 3000 571524 3012
rect 571576 3000 571582 3052
rect 194468 2944 196388 2972
rect 194468 2932 194474 2944
rect 199102 2932 199108 2984
rect 199160 2972 199166 2984
rect 204990 2972 204996 2984
rect 199160 2944 204996 2972
rect 199160 2932 199166 2944
rect 204990 2932 204996 2944
rect 205048 2932 205054 2984
rect 206922 2972 206928 2984
rect 205100 2944 206928 2972
rect 182910 2904 182916 2916
rect 177776 2876 182916 2904
rect 182910 2864 182916 2876
rect 182968 2864 182974 2916
rect 183738 2864 183744 2916
rect 183796 2904 183802 2916
rect 190638 2904 190644 2916
rect 183796 2876 190644 2904
rect 183796 2864 183802 2876
rect 190638 2864 190644 2876
rect 190696 2864 190702 2916
rect 192386 2864 192392 2916
rect 192444 2904 192450 2916
rect 198366 2904 198372 2916
rect 192444 2876 198372 2904
rect 192444 2864 192450 2876
rect 198366 2864 198372 2876
rect 198424 2864 198430 2916
rect 201494 2864 201500 2916
rect 201552 2904 201558 2916
rect 205100 2904 205128 2944
rect 206922 2932 206928 2944
rect 206980 2932 206986 2984
rect 208578 2932 208584 2984
rect 208636 2972 208642 2984
rect 213822 2972 213828 2984
rect 208636 2944 213828 2972
rect 208636 2932 208642 2944
rect 213822 2932 213828 2944
rect 213880 2932 213886 2984
rect 214466 2932 214472 2984
rect 214524 2972 214530 2984
rect 219342 2972 219348 2984
rect 214524 2944 219348 2972
rect 214524 2932 214530 2944
rect 219342 2932 219348 2944
rect 219400 2932 219406 2984
rect 223942 2932 223948 2984
rect 224000 2932 224006 2984
rect 225138 2932 225144 2984
rect 225196 2972 225202 2984
rect 229554 2972 229560 2984
rect 225196 2944 229560 2972
rect 225196 2932 225202 2944
rect 229554 2932 229560 2944
rect 229612 2932 229618 2984
rect 231026 2932 231032 2984
rect 231084 2972 231090 2984
rect 235074 2972 235080 2984
rect 231084 2944 235080 2972
rect 231084 2932 231090 2944
rect 235074 2932 235080 2944
rect 235132 2932 235138 2984
rect 235810 2932 235816 2984
rect 235868 2972 235874 2984
rect 239490 2972 239496 2984
rect 235868 2944 239496 2972
rect 235868 2932 235874 2944
rect 239490 2932 239496 2944
rect 239548 2932 239554 2984
rect 242066 2932 242072 2984
rect 242124 2972 242130 2984
rect 245010 2972 245016 2984
rect 242124 2944 245016 2972
rect 242124 2932 242130 2944
rect 245010 2932 245016 2944
rect 245068 2932 245074 2984
rect 247586 2932 247592 2984
rect 247644 2972 247650 2984
rect 250530 2972 250536 2984
rect 247644 2944 250536 2972
rect 247644 2932 247650 2944
rect 250530 2932 250536 2944
rect 250588 2932 250594 2984
rect 253474 2932 253480 2984
rect 253532 2972 253538 2984
rect 256050 2972 256056 2984
rect 253532 2944 256056 2972
rect 253532 2932 253538 2944
rect 256050 2932 256056 2944
rect 256108 2932 256114 2984
rect 310238 2932 310244 2984
rect 310296 2972 310302 2984
rect 311434 2972 311440 2984
rect 310296 2944 311440 2972
rect 310296 2932 310302 2944
rect 311434 2932 311440 2944
rect 311492 2932 311498 2984
rect 325694 2932 325700 2984
rect 325752 2972 325758 2984
rect 327994 2972 328000 2984
rect 325752 2944 328000 2972
rect 325752 2932 325758 2944
rect 327994 2932 328000 2944
rect 328052 2932 328058 2984
rect 329006 2932 329012 2984
rect 329064 2972 329070 2984
rect 331582 2972 331588 2984
rect 329064 2944 331588 2972
rect 329064 2932 329070 2944
rect 331582 2932 331588 2944
rect 331640 2932 331646 2984
rect 332318 2932 332324 2984
rect 332376 2972 332382 2984
rect 335078 2972 335084 2984
rect 332376 2944 335084 2972
rect 332376 2932 332382 2944
rect 335078 2932 335084 2944
rect 335136 2932 335142 2984
rect 341150 2932 341156 2984
rect 341208 2972 341214 2984
rect 344554 2972 344560 2984
rect 341208 2944 344560 2972
rect 341208 2932 341214 2944
rect 344554 2932 344560 2944
rect 344612 2932 344618 2984
rect 513282 2932 513288 2984
rect 513340 2972 513346 2984
rect 529014 2972 529020 2984
rect 513340 2944 529020 2972
rect 513340 2932 513346 2944
rect 529014 2932 529020 2944
rect 529072 2932 529078 2984
rect 549806 2932 549812 2984
rect 549864 2972 549870 2984
rect 568022 2972 568028 2984
rect 549864 2944 568028 2972
rect 549864 2932 549870 2944
rect 568022 2932 568028 2944
rect 568080 2932 568086 2984
rect 201552 2876 205128 2904
rect 201552 2864 201558 2876
rect 206186 2864 206192 2916
rect 206244 2904 206250 2916
rect 211614 2904 211620 2916
rect 206244 2876 211620 2904
rect 206244 2864 206250 2876
rect 211614 2864 211620 2876
rect 211672 2864 211678 2916
rect 213362 2864 213368 2916
rect 213420 2904 213426 2916
rect 217962 2904 217968 2916
rect 213420 2876 217968 2904
rect 213420 2864 213426 2876
rect 217962 2864 217968 2876
rect 218020 2864 218026 2916
rect 218054 2864 218060 2916
rect 218112 2904 218118 2916
rect 222930 2904 222936 2916
rect 218112 2876 222936 2904
rect 218112 2864 218118 2876
rect 222930 2864 222936 2876
rect 222988 2864 222994 2916
rect 223114 2864 223120 2916
rect 223172 2904 223178 2916
rect 227346 2904 227352 2916
rect 223172 2876 227352 2904
rect 223172 2864 223178 2876
rect 227346 2864 227352 2876
rect 227404 2864 227410 2916
rect 227530 2864 227536 2916
rect 227588 2904 227594 2916
rect 231762 2904 231768 2916
rect 227588 2876 231768 2904
rect 227588 2864 227594 2876
rect 231762 2864 231768 2876
rect 231820 2864 231826 2916
rect 232222 2864 232228 2916
rect 232280 2904 232286 2916
rect 236178 2904 236184 2916
rect 232280 2876 236184 2904
rect 232280 2864 232286 2876
rect 236178 2864 236184 2876
rect 236236 2864 236242 2916
rect 237006 2864 237012 2916
rect 237064 2904 237070 2916
rect 240594 2904 240600 2916
rect 237064 2876 240600 2904
rect 237064 2864 237070 2876
rect 240594 2864 240600 2876
rect 240652 2864 240658 2916
rect 244090 2864 244096 2916
rect 244148 2904 244154 2916
rect 247218 2904 247224 2916
rect 244148 2876 247224 2904
rect 244148 2864 244154 2876
rect 247218 2864 247224 2876
rect 247276 2864 247282 2916
rect 249978 2864 249984 2916
rect 250036 2904 250042 2916
rect 252738 2904 252744 2916
rect 250036 2876 252744 2904
rect 250036 2864 250042 2876
rect 252738 2864 252744 2876
rect 252796 2864 252802 2916
rect 254670 2864 254676 2916
rect 254728 2904 254734 2916
rect 257154 2904 257160 2916
rect 254728 2876 257160 2904
rect 254728 2864 254734 2876
rect 257154 2864 257160 2876
rect 257212 2864 257218 2916
rect 261754 2864 261760 2916
rect 261812 2904 261818 2916
rect 263778 2904 263784 2916
rect 261812 2876 263784 2904
rect 261812 2864 261818 2876
rect 263778 2864 263784 2876
rect 263836 2864 263842 2916
rect 312446 2864 312452 2916
rect 312504 2904 312510 2916
rect 313826 2904 313832 2916
rect 312504 2876 313832 2904
rect 312504 2864 312510 2876
rect 313826 2864 313832 2876
rect 313884 2864 313890 2916
rect 314562 2864 314568 2916
rect 314620 2904 314626 2916
rect 316218 2904 316224 2916
rect 314620 2876 316224 2904
rect 314620 2864 314626 2876
rect 316218 2864 316224 2876
rect 316276 2864 316282 2916
rect 316862 2864 316868 2916
rect 316920 2904 316926 2916
rect 318518 2904 318524 2916
rect 316920 2876 318524 2904
rect 316920 2864 316926 2876
rect 318518 2864 318524 2876
rect 318576 2864 318582 2916
rect 319070 2864 319076 2916
rect 319128 2904 319134 2916
rect 320910 2904 320916 2916
rect 319128 2876 320916 2904
rect 319128 2864 319134 2876
rect 320910 2864 320916 2876
rect 320968 2864 320974 2916
rect 321278 2864 321284 2916
rect 321336 2904 321342 2916
rect 323302 2904 323308 2916
rect 321336 2876 323308 2904
rect 321336 2864 321342 2876
rect 323302 2864 323308 2876
rect 323360 2864 323366 2916
rect 323486 2864 323492 2916
rect 323544 2904 323550 2916
rect 325602 2904 325608 2916
rect 323544 2876 325608 2904
rect 323544 2864 323550 2876
rect 325602 2864 325608 2876
rect 325660 2864 325666 2916
rect 327902 2864 327908 2916
rect 327960 2904 327966 2916
rect 330386 2904 330392 2916
rect 327960 2876 330392 2904
rect 327960 2864 327966 2876
rect 330386 2864 330392 2876
rect 330444 2864 330450 2916
rect 331122 2864 331128 2916
rect 331180 2904 331186 2916
rect 333882 2904 333888 2916
rect 331180 2876 333888 2904
rect 331180 2864 331186 2876
rect 333882 2864 333888 2876
rect 333940 2864 333946 2916
rect 334526 2864 334532 2916
rect 334584 2904 334590 2916
rect 337470 2904 337476 2916
rect 334584 2876 337476 2904
rect 334584 2864 334590 2876
rect 337470 2864 337476 2876
rect 337528 2864 337534 2916
rect 340046 2864 340052 2916
rect 340104 2904 340110 2916
rect 342990 2904 342996 2916
rect 340104 2876 342996 2904
rect 340104 2864 340110 2876
rect 342990 2864 342996 2876
rect 343048 2864 343054 2916
rect 517514 2864 517520 2916
rect 517572 2904 517578 2916
rect 523034 2904 523040 2916
rect 517572 2876 523040 2904
rect 517572 2864 517578 2876
rect 523034 2864 523040 2876
rect 523092 2864 523098 2916
rect 525794 2864 525800 2916
rect 525852 2904 525858 2916
rect 531314 2904 531320 2916
rect 525852 2876 531320 2904
rect 525852 2864 525858 2876
rect 531314 2864 531320 2876
rect 531372 2864 531378 2916
rect 536558 2864 536564 2916
rect 536616 2904 536622 2916
rect 553762 2904 553768 2916
rect 536616 2876 553768 2904
rect 536616 2864 536622 2876
rect 553762 2864 553768 2876
rect 553820 2864 553826 2916
rect 559742 2864 559748 2916
rect 559800 2904 559806 2916
rect 578602 2904 578608 2916
rect 559800 2876 578608 2904
rect 559800 2864 559806 2876
rect 578602 2864 578608 2876
rect 578660 2864 578666 2916
rect 154206 2836 154212 2848
rect 147646 2808 154212 2836
rect 154206 2796 154212 2808
rect 154264 2796 154270 2848
rect 158898 2796 158904 2848
rect 158956 2836 158962 2848
rect 167730 2836 167736 2848
rect 158956 2808 167736 2836
rect 158956 2796 158962 2808
rect 167730 2796 167736 2808
rect 167788 2796 167794 2848
rect 168374 2796 168380 2848
rect 168432 2836 168438 2848
rect 176286 2836 176292 2848
rect 168432 2808 176292 2836
rect 168432 2796 168438 2808
rect 176286 2796 176292 2808
rect 176344 2796 176350 2848
rect 180242 2796 180248 2848
rect 180300 2836 180306 2848
rect 187326 2836 187332 2848
rect 180300 2808 187332 2836
rect 180300 2796 180306 2808
rect 187326 2796 187332 2808
rect 187384 2796 187390 2848
rect 199470 2836 199476 2848
rect 193232 2808 199476 2836
rect 193232 2780 193260 2808
rect 199470 2796 199476 2808
rect 199528 2796 199534 2848
rect 205082 2796 205088 2848
rect 205140 2836 205146 2848
rect 210510 2836 210516 2848
rect 205140 2808 210516 2836
rect 205140 2796 205146 2808
rect 210510 2796 210516 2808
rect 210568 2796 210574 2848
rect 210970 2796 210976 2848
rect 211028 2836 211034 2848
rect 216030 2836 216036 2848
rect 211028 2808 216036 2836
rect 211028 2796 211034 2808
rect 216030 2796 216036 2808
rect 216088 2796 216094 2848
rect 216858 2796 216864 2848
rect 216916 2836 216922 2848
rect 221826 2836 221832 2848
rect 216916 2808 221832 2836
rect 216916 2796 216922 2808
rect 221826 2796 221832 2808
rect 221884 2796 221890 2848
rect 226334 2796 226340 2848
rect 226392 2836 226398 2848
rect 230658 2836 230664 2848
rect 226392 2808 230664 2836
rect 226392 2796 226398 2808
rect 230658 2796 230664 2808
rect 230716 2796 230722 2848
rect 233418 2796 233424 2848
rect 233476 2836 233482 2848
rect 237282 2836 237288 2848
rect 233476 2808 237288 2836
rect 233476 2796 233482 2808
rect 237282 2796 237288 2808
rect 237340 2796 237346 2848
rect 238110 2796 238116 2848
rect 238168 2836 238174 2848
rect 241698 2836 241704 2848
rect 238168 2808 241704 2836
rect 238168 2796 238174 2808
rect 241698 2796 241704 2808
rect 241756 2796 241762 2848
rect 242894 2796 242900 2848
rect 242952 2836 242958 2848
rect 246114 2836 246120 2848
rect 242952 2808 246120 2836
rect 242952 2796 242958 2808
rect 246114 2796 246120 2808
rect 246172 2796 246178 2848
rect 246390 2796 246396 2848
rect 246448 2836 246454 2848
rect 249426 2836 249432 2848
rect 246448 2808 249432 2836
rect 246448 2796 246454 2808
rect 249426 2796 249432 2808
rect 249484 2796 249490 2848
rect 252370 2796 252376 2848
rect 252428 2836 252434 2848
rect 254946 2836 254952 2848
rect 252428 2808 254952 2836
rect 252428 2796 252434 2808
rect 254946 2796 254952 2808
rect 255004 2796 255010 2848
rect 255866 2796 255872 2848
rect 255924 2836 255930 2848
rect 258258 2836 258264 2848
rect 255924 2808 258264 2836
rect 255924 2796 255930 2808
rect 258258 2796 258264 2808
rect 258316 2796 258322 2848
rect 260650 2796 260656 2848
rect 260708 2836 260714 2848
rect 262674 2836 262680 2848
rect 260708 2808 262680 2836
rect 260708 2796 260714 2808
rect 262674 2796 262680 2808
rect 262732 2796 262738 2848
rect 304718 2796 304724 2848
rect 304776 2836 304782 2848
rect 305546 2836 305552 2848
rect 304776 2808 305552 2836
rect 304776 2796 304782 2808
rect 305546 2796 305552 2808
rect 305604 2796 305610 2848
rect 306926 2796 306932 2848
rect 306984 2836 306990 2848
rect 307938 2836 307944 2848
rect 306984 2808 307944 2836
rect 306984 2796 306990 2808
rect 307938 2796 307944 2808
rect 307996 2796 308002 2848
rect 309134 2796 309140 2848
rect 309192 2836 309198 2848
rect 310238 2836 310244 2848
rect 309192 2808 310244 2836
rect 309192 2796 309198 2808
rect 310238 2796 310244 2808
rect 310296 2796 310302 2848
rect 311342 2796 311348 2848
rect 311400 2836 311406 2848
rect 312630 2836 312636 2848
rect 311400 2808 312636 2836
rect 311400 2796 311406 2808
rect 312630 2796 312636 2808
rect 312688 2796 312694 2848
rect 313550 2796 313556 2848
rect 313608 2836 313614 2848
rect 315022 2836 315028 2848
rect 313608 2808 315028 2836
rect 313608 2796 313614 2808
rect 315022 2796 315028 2808
rect 315080 2796 315086 2848
rect 315758 2796 315764 2848
rect 315816 2836 315822 2848
rect 317322 2836 317328 2848
rect 315816 2808 317328 2836
rect 315816 2796 315822 2808
rect 317322 2796 317328 2808
rect 317380 2796 317386 2848
rect 317966 2796 317972 2848
rect 318024 2836 318030 2848
rect 319714 2836 319720 2848
rect 318024 2808 319720 2836
rect 318024 2796 318030 2808
rect 319714 2796 319720 2808
rect 319772 2796 319778 2848
rect 320082 2796 320088 2848
rect 320140 2836 320146 2848
rect 322106 2836 322112 2848
rect 320140 2808 322112 2836
rect 320140 2796 320146 2808
rect 322106 2796 322112 2808
rect 322164 2796 322170 2848
rect 322382 2796 322388 2848
rect 322440 2836 322446 2848
rect 324406 2836 324412 2848
rect 322440 2808 324412 2836
rect 322440 2796 322446 2808
rect 324406 2796 324412 2808
rect 324464 2796 324470 2848
rect 324590 2796 324596 2848
rect 324648 2836 324654 2848
rect 326798 2836 326804 2848
rect 324648 2808 326804 2836
rect 324648 2796 324654 2808
rect 326798 2796 326804 2808
rect 326856 2796 326862 2848
rect 326982 2796 326988 2848
rect 327040 2836 327046 2848
rect 329190 2836 329196 2848
rect 327040 2808 329196 2836
rect 327040 2796 327046 2808
rect 329190 2796 329196 2808
rect 329248 2796 329254 2848
rect 330110 2796 330116 2848
rect 330168 2836 330174 2848
rect 332686 2836 332692 2848
rect 330168 2808 332692 2836
rect 330168 2796 330174 2808
rect 332686 2796 332692 2808
rect 332744 2796 332750 2848
rect 335630 2796 335636 2848
rect 335688 2836 335694 2848
rect 338666 2836 338672 2848
rect 335688 2808 338672 2836
rect 335688 2796 335694 2808
rect 338666 2796 338672 2808
rect 338724 2796 338730 2848
rect 338942 2796 338948 2848
rect 339000 2836 339006 2848
rect 342070 2836 342076 2848
rect 339000 2808 342076 2836
rect 339000 2796 339006 2808
rect 342070 2796 342076 2808
rect 342128 2796 342134 2848
rect 346670 2796 346676 2848
rect 346728 2836 346734 2848
rect 350442 2836 350448 2848
rect 346728 2808 350448 2836
rect 346728 2796 346734 2808
rect 350442 2796 350448 2808
rect 350500 2796 350506 2848
rect 353202 2796 353208 2848
rect 353260 2836 353266 2848
rect 357526 2836 357532 2848
rect 353260 2808 357532 2836
rect 353260 2796 353266 2808
rect 357526 2796 357532 2808
rect 357584 2796 357590 2848
rect 372338 2796 372344 2848
rect 372396 2836 372402 2848
rect 377674 2836 377680 2848
rect 372396 2808 377680 2836
rect 372396 2796 372402 2808
rect 377674 2796 377680 2808
rect 377732 2796 377738 2848
rect 517606 2796 517612 2848
rect 517664 2836 517670 2848
rect 521838 2836 521844 2848
rect 517664 2808 521844 2836
rect 517664 2796 517670 2808
rect 521838 2796 521844 2808
rect 521896 2796 521902 2848
rect 562962 2796 562968 2848
rect 563020 2836 563026 2848
rect 582190 2836 582196 2848
rect 563020 2808 582196 2836
rect 563020 2796 563026 2808
rect 582190 2796 582196 2808
rect 582248 2796 582254 2848
rect 193214 2728 193220 2780
rect 193272 2728 193278 2780
rect 176654 1300 176660 1352
rect 176712 1340 176718 1352
rect 184290 1340 184296 1352
rect 176712 1312 184296 1340
rect 176712 1300 176718 1312
rect 184290 1300 184296 1312
rect 184348 1300 184354 1352
rect 187326 1300 187332 1352
rect 187384 1340 187390 1352
rect 194226 1340 194232 1352
rect 187384 1312 194232 1340
rect 187384 1300 187390 1312
rect 194226 1300 194232 1312
rect 194284 1300 194290 1352
rect 198274 1300 198280 1352
rect 198332 1340 198338 1352
rect 204162 1340 204168 1352
rect 198332 1312 204168 1340
rect 198332 1300 198338 1312
rect 204162 1300 204168 1312
rect 204220 1300 204226 1352
rect 207382 1300 207388 1352
rect 207440 1340 207446 1352
rect 212994 1340 213000 1352
rect 207440 1312 213000 1340
rect 207440 1300 207446 1312
rect 212994 1300 213000 1312
rect 213052 1300 213058 1352
rect 257062 1300 257068 1352
rect 257120 1340 257126 1352
rect 259362 1340 259368 1352
rect 257120 1312 259368 1340
rect 257120 1300 257126 1312
rect 259362 1300 259368 1312
rect 259420 1300 259426 1352
rect 259454 1300 259460 1352
rect 259512 1340 259518 1352
rect 261570 1340 261576 1352
rect 259512 1312 261576 1340
rect 259512 1300 259518 1312
rect 261570 1300 261576 1312
rect 261628 1300 261634 1352
rect 262950 1300 262956 1352
rect 263008 1340 263014 1352
rect 264882 1340 264888 1352
rect 263008 1312 264888 1340
rect 263008 1300 263014 1312
rect 264882 1300 264888 1312
rect 264940 1300 264946 1352
rect 265342 1300 265348 1352
rect 265400 1340 265406 1352
rect 267090 1340 267096 1352
rect 265400 1312 267096 1340
rect 265400 1300 265406 1312
rect 267090 1300 267096 1312
rect 267148 1300 267154 1352
rect 267734 1300 267740 1352
rect 267792 1340 267798 1352
rect 269298 1340 269304 1352
rect 267792 1312 269304 1340
rect 267792 1300 267798 1312
rect 269298 1300 269304 1312
rect 269356 1300 269362 1352
rect 271230 1300 271236 1352
rect 271288 1340 271294 1352
rect 272610 1340 272616 1352
rect 271288 1312 272616 1340
rect 271288 1300 271294 1312
rect 272610 1300 272616 1312
rect 272668 1300 272674 1352
rect 273622 1300 273628 1352
rect 273680 1340 273686 1352
rect 274818 1340 274824 1352
rect 273680 1312 274824 1340
rect 273680 1300 273686 1312
rect 274818 1300 274824 1312
rect 274876 1300 274882 1352
rect 277118 1300 277124 1352
rect 277176 1340 277182 1352
rect 278130 1340 278136 1352
rect 277176 1312 278136 1340
rect 277176 1300 277182 1312
rect 278130 1300 278136 1312
rect 278188 1300 278194 1352
rect 279510 1300 279516 1352
rect 279568 1340 279574 1352
rect 280338 1340 280344 1352
rect 279568 1312 280344 1340
rect 279568 1300 279574 1312
rect 280338 1300 280344 1312
rect 280396 1300 280402 1352
rect 336642 1300 336648 1352
rect 336700 1340 336706 1352
rect 339862 1340 339868 1352
rect 336700 1312 339868 1340
rect 336700 1300 336706 1312
rect 339862 1300 339868 1312
rect 339920 1300 339926 1352
rect 342162 1300 342168 1352
rect 342220 1340 342226 1352
rect 345750 1340 345756 1352
rect 342220 1312 345756 1340
rect 342220 1300 342226 1312
rect 345750 1300 345756 1312
rect 345808 1300 345814 1352
rect 348878 1300 348884 1352
rect 348936 1340 348942 1352
rect 352834 1340 352840 1352
rect 348936 1312 352840 1340
rect 348936 1300 348942 1312
rect 352834 1300 352840 1312
rect 352892 1300 352898 1352
rect 356606 1300 356612 1352
rect 356664 1340 356670 1352
rect 361114 1340 361120 1352
rect 356664 1312 361120 1340
rect 356664 1300 356670 1312
rect 361114 1300 361120 1312
rect 361172 1300 361178 1352
rect 364242 1300 364248 1352
rect 364300 1340 364306 1352
rect 369394 1340 369400 1352
rect 364300 1312 369400 1340
rect 364300 1300 364306 1312
rect 369394 1300 369400 1312
rect 369452 1300 369458 1352
rect 374270 1300 374276 1352
rect 374328 1340 374334 1352
rect 379606 1340 379612 1352
rect 374328 1312 379612 1340
rect 374328 1300 374334 1312
rect 379606 1300 379612 1312
rect 379664 1300 379670 1352
rect 384206 1300 384212 1352
rect 384264 1340 384270 1352
rect 390646 1340 390652 1352
rect 384264 1312 390652 1340
rect 384264 1300 384270 1312
rect 390646 1300 390652 1312
rect 390704 1300 390710 1352
rect 396350 1300 396356 1352
rect 396408 1340 396414 1352
rect 403618 1340 403624 1352
rect 396408 1312 403624 1340
rect 396408 1300 396414 1312
rect 403618 1300 403624 1312
rect 403676 1300 403682 1352
rect 406286 1300 406292 1352
rect 406344 1340 406350 1352
rect 414290 1340 414296 1352
rect 406344 1312 414296 1340
rect 406344 1300 406350 1312
rect 414290 1300 414296 1312
rect 414348 1300 414354 1352
rect 419442 1300 419448 1352
rect 419500 1340 419506 1352
rect 428274 1340 428280 1352
rect 419500 1312 428280 1340
rect 419500 1300 419506 1312
rect 428274 1300 428280 1312
rect 428332 1300 428338 1352
rect 428366 1300 428372 1352
rect 428424 1340 428430 1352
rect 428424 1312 435956 1340
rect 428424 1300 428430 1312
rect 98638 1232 98644 1284
rect 98696 1272 98702 1284
rect 105906 1272 105912 1284
rect 98696 1244 105912 1272
rect 98696 1232 98702 1244
rect 105906 1232 105912 1244
rect 105964 1232 105970 1284
rect 188890 1232 188896 1284
rect 188948 1272 188954 1284
rect 195330 1272 195336 1284
rect 188948 1244 195336 1272
rect 188948 1232 188954 1244
rect 195330 1232 195336 1244
rect 195388 1232 195394 1284
rect 197170 1232 197176 1284
rect 197228 1272 197234 1284
rect 203058 1272 203064 1284
rect 197228 1244 203064 1272
rect 197228 1232 197234 1244
rect 203058 1232 203064 1244
rect 203116 1232 203122 1284
rect 258258 1232 258264 1284
rect 258316 1272 258322 1284
rect 260466 1272 260472 1284
rect 258316 1244 260472 1272
rect 258316 1232 258322 1244
rect 260466 1232 260472 1244
rect 260524 1232 260530 1284
rect 264146 1232 264152 1284
rect 264204 1272 264210 1284
rect 265986 1272 265992 1284
rect 264204 1244 265992 1272
rect 264204 1232 264210 1244
rect 265986 1232 265992 1244
rect 266044 1232 266050 1284
rect 266538 1232 266544 1284
rect 266596 1272 266602 1284
rect 268194 1272 268200 1284
rect 266596 1244 268200 1272
rect 266596 1232 266602 1244
rect 268194 1232 268200 1244
rect 268252 1232 268258 1284
rect 270034 1232 270040 1284
rect 270092 1272 270098 1284
rect 271506 1272 271512 1284
rect 270092 1244 271512 1272
rect 270092 1232 270098 1244
rect 271506 1232 271512 1244
rect 271564 1232 271570 1284
rect 272426 1232 272432 1284
rect 272484 1272 272490 1284
rect 273714 1272 273720 1284
rect 272484 1244 273720 1272
rect 272484 1232 272490 1244
rect 273714 1232 273720 1244
rect 273772 1232 273778 1284
rect 343358 1232 343364 1284
rect 343416 1272 343422 1284
rect 346946 1272 346952 1284
rect 343416 1244 346952 1272
rect 343416 1232 343422 1244
rect 346946 1232 346952 1244
rect 347004 1232 347010 1284
rect 349982 1232 349988 1284
rect 350040 1272 350046 1284
rect 354030 1272 354036 1284
rect 350040 1244 354036 1272
rect 350040 1232 350046 1244
rect 354030 1232 354036 1244
rect 354088 1232 354094 1284
rect 357710 1232 357716 1284
rect 357768 1272 357774 1284
rect 362310 1272 362316 1284
rect 357768 1244 362316 1272
rect 357768 1232 357774 1244
rect 362310 1232 362316 1244
rect 362368 1232 362374 1284
rect 365438 1232 365444 1284
rect 365496 1272 365502 1284
rect 370222 1272 370228 1284
rect 365496 1244 370228 1272
rect 365496 1232 365502 1244
rect 370222 1232 370228 1244
rect 370280 1232 370286 1284
rect 370958 1232 370964 1284
rect 371016 1272 371022 1284
rect 376110 1272 376116 1284
rect 371016 1244 376116 1272
rect 371016 1232 371022 1244
rect 376110 1232 376116 1244
rect 376168 1232 376174 1284
rect 377582 1232 377588 1284
rect 377640 1272 377646 1284
rect 383562 1272 383568 1284
rect 377640 1244 383568 1272
rect 377640 1232 377646 1244
rect 383562 1232 383568 1244
rect 383620 1232 383626 1284
rect 388622 1232 388628 1284
rect 388680 1272 388686 1284
rect 395338 1272 395344 1284
rect 388680 1244 395344 1272
rect 388680 1232 388686 1244
rect 395338 1232 395344 1244
rect 395396 1232 395402 1284
rect 404078 1232 404084 1284
rect 404136 1272 404142 1284
rect 411898 1272 411904 1284
rect 404136 1244 411904 1272
rect 404136 1232 404142 1244
rect 411898 1232 411904 1244
rect 411956 1232 411962 1284
rect 413922 1232 413928 1284
rect 413980 1272 413986 1284
rect 422570 1272 422576 1284
rect 413980 1244 422576 1272
rect 413980 1232 413986 1244
rect 422570 1232 422576 1244
rect 422628 1232 422634 1284
rect 426158 1232 426164 1284
rect 426216 1272 426222 1284
rect 435174 1272 435180 1284
rect 426216 1244 435180 1272
rect 426216 1232 426222 1244
rect 435174 1232 435180 1244
rect 435232 1232 435238 1284
rect 435928 1272 435956 1312
rect 436002 1300 436008 1352
rect 436060 1340 436066 1352
rect 436060 1312 443776 1340
rect 436060 1300 436066 1312
rect 437566 1272 437572 1284
rect 435928 1244 437572 1272
rect 437566 1232 437572 1244
rect 437624 1232 437630 1284
rect 438302 1232 438308 1284
rect 438360 1272 438366 1284
rect 443748 1272 443776 1312
rect 443822 1300 443828 1352
rect 443880 1340 443886 1352
rect 454126 1340 454132 1352
rect 443880 1312 454132 1340
rect 443880 1300 443886 1312
rect 454126 1300 454132 1312
rect 454184 1300 454190 1352
rect 456978 1340 456984 1352
rect 454788 1312 456984 1340
rect 445846 1272 445852 1284
rect 438360 1244 443684 1272
rect 443748 1244 445852 1272
rect 438360 1232 438366 1244
rect 186130 1164 186136 1216
rect 186188 1204 186194 1216
rect 193122 1204 193128 1216
rect 186188 1176 193128 1204
rect 186188 1164 186194 1176
rect 193122 1164 193128 1176
rect 193180 1164 193186 1216
rect 268838 1164 268844 1216
rect 268896 1204 268902 1216
rect 270402 1204 270408 1216
rect 268896 1176 270408 1204
rect 268896 1164 268902 1176
rect 270402 1164 270408 1176
rect 270460 1164 270466 1216
rect 359918 1164 359924 1216
rect 359976 1204 359982 1216
rect 364610 1204 364616 1216
rect 359976 1176 364616 1204
rect 359976 1164 359982 1176
rect 364610 1164 364616 1176
rect 364668 1164 364674 1216
rect 366542 1164 366548 1216
rect 366600 1204 366606 1216
rect 371326 1204 371332 1216
rect 366600 1176 371332 1204
rect 366600 1164 366606 1176
rect 371326 1164 371332 1176
rect 371384 1164 371390 1216
rect 378686 1164 378692 1216
rect 378744 1204 378750 1216
rect 384390 1204 384396 1216
rect 378744 1176 384396 1204
rect 378744 1164 378750 1176
rect 384390 1164 384396 1176
rect 384448 1164 384454 1216
rect 387518 1164 387524 1216
rect 387576 1204 387582 1216
rect 394234 1204 394240 1216
rect 387576 1176 394240 1204
rect 387576 1164 387582 1176
rect 394234 1164 394240 1176
rect 394292 1164 394298 1216
rect 395246 1164 395252 1216
rect 395304 1204 395310 1216
rect 402514 1204 402520 1216
rect 395304 1176 402520 1204
rect 395304 1164 395310 1176
rect 402514 1164 402520 1176
rect 402572 1164 402578 1216
rect 412910 1164 412916 1216
rect 412968 1204 412974 1216
rect 421374 1204 421380 1216
rect 412968 1176 421380 1204
rect 412968 1164 412974 1176
rect 421374 1164 421380 1176
rect 421432 1164 421438 1216
rect 421742 1164 421748 1216
rect 421800 1204 421806 1216
rect 430850 1204 430856 1216
rect 421800 1176 430856 1204
rect 421800 1164 421806 1176
rect 430850 1164 430856 1176
rect 430908 1164 430914 1216
rect 439406 1164 439412 1216
rect 439464 1204 439470 1216
rect 443546 1204 443552 1216
rect 439464 1176 443552 1204
rect 439464 1164 439470 1176
rect 443546 1164 443552 1176
rect 443604 1164 443610 1216
rect 443656 1204 443684 1244
rect 445846 1232 445852 1244
rect 445904 1232 445910 1284
rect 449342 1232 449348 1284
rect 449400 1272 449406 1284
rect 454788 1272 454816 1312
rect 456978 1300 456984 1312
rect 457036 1300 457042 1352
rect 457070 1300 457076 1352
rect 457128 1340 457134 1352
rect 468294 1340 468300 1352
rect 457128 1312 468300 1340
rect 457128 1300 457134 1312
rect 468294 1300 468300 1312
rect 468352 1300 468358 1352
rect 481358 1300 481364 1352
rect 481416 1340 481422 1352
rect 494698 1340 494704 1352
rect 481416 1312 494704 1340
rect 481416 1300 481422 1312
rect 494698 1300 494704 1312
rect 494756 1300 494762 1352
rect 495710 1300 495716 1352
rect 495768 1340 495774 1352
rect 509694 1340 509700 1352
rect 495768 1312 509700 1340
rect 495768 1300 495774 1312
rect 509694 1300 509700 1312
rect 509752 1300 509758 1352
rect 510062 1300 510068 1352
rect 510120 1340 510126 1352
rect 525426 1340 525432 1352
rect 510120 1312 525432 1340
rect 510120 1300 510126 1312
rect 525426 1300 525432 1312
rect 525484 1300 525490 1352
rect 539870 1300 539876 1352
rect 539928 1340 539934 1352
rect 556982 1340 556988 1352
rect 539928 1312 556988 1340
rect 539928 1300 539934 1312
rect 556982 1300 556988 1312
rect 557040 1300 557046 1352
rect 449400 1244 454816 1272
rect 449400 1232 449406 1244
rect 454862 1232 454868 1284
rect 454920 1272 454926 1284
rect 454920 1244 460934 1272
rect 454920 1232 454926 1244
rect 448606 1204 448612 1216
rect 443656 1176 448612 1204
rect 448606 1164 448612 1176
rect 448664 1164 448670 1216
rect 450446 1164 450452 1216
rect 450504 1204 450510 1216
rect 460906 1204 460934 1244
rect 462590 1232 462596 1284
rect 462648 1272 462654 1284
rect 474182 1272 474188 1284
rect 462648 1244 474188 1272
rect 462648 1232 462654 1244
rect 474182 1232 474188 1244
rect 474240 1232 474246 1284
rect 480162 1232 480168 1284
rect 480220 1272 480226 1284
rect 493134 1272 493140 1284
rect 480220 1244 493140 1272
rect 480220 1232 480226 1244
rect 493134 1232 493140 1244
rect 493192 1232 493198 1284
rect 493502 1232 493508 1284
rect 493560 1272 493566 1284
rect 507302 1272 507308 1284
rect 493560 1244 507308 1272
rect 493560 1232 493566 1244
rect 507302 1232 507308 1244
rect 507360 1232 507366 1284
rect 507762 1232 507768 1284
rect 507820 1272 507826 1284
rect 517514 1272 517520 1284
rect 507820 1244 517520 1272
rect 507820 1232 507826 1244
rect 517514 1232 517520 1244
rect 517572 1232 517578 1284
rect 534350 1232 534356 1284
rect 534408 1272 534414 1284
rect 551094 1272 551100 1284
rect 534408 1244 551100 1272
rect 534408 1232 534414 1244
rect 551094 1232 551100 1244
rect 551152 1232 551158 1284
rect 465902 1204 465908 1216
rect 450504 1176 456104 1204
rect 460906 1176 465908 1204
rect 450504 1164 450510 1176
rect 352190 1096 352196 1148
rect 352248 1136 352254 1148
rect 356330 1136 356336 1148
rect 352248 1108 356336 1136
rect 352248 1096 352254 1108
rect 356330 1096 356336 1108
rect 356388 1096 356394 1148
rect 361022 1096 361028 1148
rect 361080 1136 361086 1148
rect 365438 1136 365444 1148
rect 361080 1108 365444 1136
rect 361080 1096 361086 1108
rect 365438 1096 365444 1108
rect 365496 1096 365502 1148
rect 367646 1096 367652 1148
rect 367704 1136 367710 1148
rect 372890 1136 372896 1148
rect 367704 1108 372896 1136
rect 367704 1096 367710 1108
rect 372890 1096 372896 1108
rect 372948 1096 372954 1148
rect 375282 1096 375288 1148
rect 375340 1136 375346 1148
rect 375340 1108 379744 1136
rect 375340 1096 375346 1108
rect 4062 1028 4068 1080
rect 4120 1068 4126 1080
rect 23106 1068 23112 1080
rect 4120 1040 23112 1068
rect 4120 1028 4126 1040
rect 23106 1028 23112 1040
rect 23164 1028 23170 1080
rect 355502 1028 355508 1080
rect 355560 1068 355566 1080
rect 359918 1068 359924 1080
rect 355560 1040 359924 1068
rect 355560 1028 355566 1040
rect 359918 1028 359924 1040
rect 359976 1028 359982 1080
rect 373166 1028 373172 1080
rect 373224 1068 373230 1080
rect 378502 1068 378508 1080
rect 373224 1040 378508 1068
rect 373224 1028 373230 1040
rect 378502 1028 378508 1040
rect 378560 1028 378566 1080
rect 379716 1068 379744 1108
rect 379790 1096 379796 1148
rect 379848 1136 379854 1148
rect 385954 1136 385960 1148
rect 379848 1108 385960 1136
rect 379848 1096 379854 1108
rect 385954 1096 385960 1108
rect 386012 1096 386018 1148
rect 386322 1096 386328 1148
rect 386380 1136 386386 1148
rect 392670 1136 392676 1148
rect 386380 1108 392676 1136
rect 386380 1096 386386 1108
rect 392670 1096 392676 1108
rect 392728 1096 392734 1148
rect 397362 1096 397368 1148
rect 397420 1136 397426 1148
rect 404814 1136 404820 1148
rect 397420 1108 404820 1136
rect 397420 1096 397426 1108
rect 404814 1096 404820 1108
rect 404872 1096 404878 1148
rect 420638 1096 420644 1148
rect 420696 1136 420702 1148
rect 429286 1136 429292 1148
rect 420696 1108 429292 1136
rect 420696 1096 420702 1108
rect 429286 1096 429292 1108
rect 429344 1096 429350 1148
rect 434990 1096 434996 1148
rect 435048 1136 435054 1148
rect 445018 1136 445024 1148
rect 435048 1108 445024 1136
rect 435048 1096 435054 1108
rect 445018 1096 445024 1108
rect 445076 1096 445082 1148
rect 445202 1096 445208 1148
rect 445260 1136 445266 1148
rect 455690 1136 455696 1148
rect 445260 1108 455696 1136
rect 445260 1096 445266 1108
rect 455690 1096 455696 1108
rect 455748 1096 455754 1148
rect 456076 1136 456104 1176
rect 465902 1164 465908 1176
rect 465960 1164 465966 1216
rect 475838 1164 475844 1216
rect 475896 1204 475902 1216
rect 488810 1204 488816 1216
rect 475896 1176 488816 1204
rect 475896 1164 475902 1176
rect 488810 1164 488816 1176
rect 488868 1164 488874 1216
rect 501230 1164 501236 1216
rect 501288 1204 501294 1216
rect 515490 1204 515496 1216
rect 501288 1176 515496 1204
rect 501288 1164 501294 1176
rect 515490 1164 515496 1176
rect 515548 1164 515554 1216
rect 516686 1164 516692 1216
rect 516744 1204 516750 1216
rect 532050 1204 532056 1216
rect 516744 1176 532056 1204
rect 516744 1164 516750 1176
rect 532050 1164 532056 1176
rect 532108 1164 532114 1216
rect 461578 1136 461584 1148
rect 456076 1108 461584 1136
rect 461578 1096 461584 1108
rect 461636 1096 461642 1148
rect 469122 1096 469128 1148
rect 469180 1136 469186 1148
rect 481358 1136 481364 1148
rect 469180 1108 481364 1136
rect 469180 1096 469186 1108
rect 481358 1096 481364 1108
rect 481416 1096 481422 1148
rect 487982 1096 487988 1148
rect 488040 1136 488046 1148
rect 501414 1136 501420 1148
rect 488040 1108 501420 1136
rect 488040 1096 488046 1108
rect 501414 1096 501420 1108
rect 501472 1096 501478 1148
rect 506750 1096 506756 1148
rect 506808 1136 506814 1148
rect 517606 1136 517612 1148
rect 506808 1108 517612 1136
rect 506808 1096 506814 1108
rect 517606 1096 517612 1108
rect 517664 1096 517670 1148
rect 522206 1096 522212 1148
rect 522264 1136 522270 1148
rect 538122 1136 538128 1148
rect 522264 1108 538128 1136
rect 522264 1096 522270 1108
rect 538122 1096 538128 1108
rect 538180 1096 538186 1148
rect 381170 1068 381176 1080
rect 379716 1040 381176 1068
rect 381170 1028 381176 1040
rect 381228 1028 381234 1080
rect 385310 1028 385316 1080
rect 385368 1068 385374 1080
rect 391842 1068 391848 1080
rect 385368 1040 391848 1068
rect 385368 1028 385374 1040
rect 391842 1028 391848 1040
rect 391900 1028 391906 1080
rect 394142 1028 394148 1080
rect 394200 1068 394206 1080
rect 401318 1068 401324 1080
rect 394200 1040 401324 1068
rect 394200 1028 394206 1040
rect 401318 1028 401324 1040
rect 401376 1028 401382 1080
rect 415118 1028 415124 1080
rect 415176 1068 415182 1080
rect 423398 1068 423404 1080
rect 415176 1040 423404 1068
rect 415176 1028 415182 1040
rect 423398 1028 423404 1040
rect 423456 1028 423462 1080
rect 424962 1028 424968 1080
rect 425020 1068 425026 1080
rect 434070 1068 434076 1080
rect 425020 1040 434076 1068
rect 425020 1028 425026 1040
rect 434070 1028 434076 1040
rect 434128 1028 434134 1080
rect 441522 1028 441528 1080
rect 441580 1068 441586 1080
rect 451734 1068 451740 1080
rect 441580 1040 451740 1068
rect 441580 1028 441586 1040
rect 451734 1028 451740 1040
rect 451792 1028 451798 1080
rect 455966 1028 455972 1080
rect 456024 1068 456030 1080
rect 467466 1068 467472 1080
rect 456024 1040 467472 1068
rect 456024 1028 456030 1040
rect 467466 1028 467472 1040
rect 467524 1028 467530 1080
rect 474642 1028 474648 1080
rect 474700 1068 474706 1080
rect 487246 1068 487252 1080
rect 474700 1040 487252 1068
rect 474700 1028 474706 1040
rect 487246 1028 487252 1040
rect 487304 1028 487310 1080
rect 518802 1028 518808 1080
rect 518860 1068 518866 1080
rect 534534 1068 534540 1080
rect 518860 1040 534540 1068
rect 518860 1028 518866 1040
rect 534534 1028 534540 1040
rect 534592 1028 534598 1080
rect 20622 960 20628 1012
rect 20680 1000 20686 1012
rect 38562 1000 38568 1012
rect 20680 972 38568 1000
rect 20680 960 20686 972
rect 38562 960 38568 972
rect 38620 960 38626 1012
rect 345566 960 345572 1012
rect 345624 1000 345630 1012
rect 349246 1000 349252 1012
rect 345624 972 349252 1000
rect 345624 960 345630 972
rect 349246 960 349252 972
rect 349304 960 349310 1012
rect 351086 960 351092 1012
rect 351144 1000 351150 1012
rect 355226 1000 355232 1012
rect 351144 972 355232 1000
rect 351144 960 351150 972
rect 355226 960 355232 972
rect 355284 960 355290 1012
rect 362126 960 362132 1012
rect 362184 1000 362190 1012
rect 367002 1000 367008 1012
rect 362184 972 367008 1000
rect 362184 960 362190 972
rect 367002 960 367008 972
rect 367060 960 367066 1012
rect 369762 960 369768 1012
rect 369820 1000 369826 1012
rect 375282 1000 375288 1012
rect 369820 972 375288 1000
rect 369820 960 369826 972
rect 375282 960 375288 972
rect 375340 960 375346 1012
rect 376478 960 376484 1012
rect 376536 1000 376542 1012
rect 382366 1000 382372 1012
rect 376536 972 382372 1000
rect 376536 960 376542 972
rect 382366 960 382372 972
rect 382424 960 382430 1012
rect 422846 960 422852 1012
rect 422904 1000 422910 1012
rect 431862 1000 431868 1012
rect 422904 972 431868 1000
rect 422904 960 422910 972
rect 431862 960 431868 972
rect 431920 960 431926 1012
rect 432782 960 432788 1012
rect 432840 1000 432846 1012
rect 442626 1000 442632 1012
rect 432840 972 442632 1000
rect 432840 960 432846 972
rect 442626 960 442632 972
rect 442684 960 442690 1012
rect 443546 960 443552 1012
rect 443604 1000 443610 1012
rect 449802 1000 449808 1012
rect 443604 972 449808 1000
rect 443604 960 443610 972
rect 449802 960 449808 972
rect 449860 960 449866 1012
rect 489086 960 489092 1012
rect 489144 1000 489150 1012
rect 502978 1000 502984 1012
rect 489144 972 502984 1000
rect 489144 960 489150 972
rect 502978 960 502984 972
rect 503036 960 503042 1012
rect 519998 960 520004 1012
rect 520056 1000 520062 1012
rect 536098 1000 536104 1012
rect 520056 972 536104 1000
rect 520056 960 520062 972
rect 536098 960 536104 972
rect 536156 960 536162 1012
rect 1670 892 1676 944
rect 1728 932 1734 944
rect 20898 932 20904 944
rect 1728 904 20904 932
rect 1728 892 1734 904
rect 20898 892 20904 904
rect 20956 892 20962 944
rect 358722 892 358728 944
rect 358780 932 358786 944
rect 363506 932 363512 944
rect 358780 904 363512 932
rect 358780 892 358786 904
rect 363506 892 363512 904
rect 363564 892 363570 944
rect 416222 892 416228 944
rect 416280 932 416286 944
rect 424962 932 424968 944
rect 416280 904 424968 932
rect 416280 892 416286 904
rect 424962 892 424968 904
rect 425020 892 425026 944
rect 433886 892 433892 944
rect 433944 932 433950 944
rect 443454 932 443460 944
rect 433944 904 443460 932
rect 433944 892 433950 904
rect 443454 892 443460 904
rect 443512 892 443518 944
rect 446030 892 446036 944
rect 446088 932 446094 944
rect 456886 932 456892 944
rect 446088 904 456892 932
rect 446088 892 446094 904
rect 456886 892 456892 904
rect 456944 892 456950 944
rect 494606 892 494612 944
rect 494664 932 494670 944
rect 508866 932 508872 944
rect 494664 904 508872 932
rect 494664 892 494670 904
rect 508866 892 508872 904
rect 508924 892 508930 944
rect 515582 892 515588 944
rect 515640 932 515646 944
rect 525794 932 525800 944
rect 515640 904 525800 932
rect 515640 892 515646 904
rect 525794 892 525800 904
rect 525852 892 525858 944
rect 532142 892 532148 944
rect 532200 932 532206 944
rect 548702 932 548708 944
rect 532200 904 548708 932
rect 532200 892 532206 904
rect 548702 892 548708 904
rect 548760 892 548766 944
rect 19426 824 19432 876
rect 19484 864 19490 876
rect 37458 864 37464 876
rect 19484 836 37464 864
rect 19484 824 19490 836
rect 37458 824 37464 836
rect 37516 824 37522 876
rect 337838 824 337844 876
rect 337896 864 337902 876
rect 340966 864 340972 876
rect 337896 836 340972 864
rect 337896 824 337902 836
rect 340966 824 340972 836
rect 341024 824 341030 876
rect 347682 824 347688 876
rect 347740 864 347746 876
rect 351638 864 351644 876
rect 347740 836 351644 864
rect 347740 824 347746 836
rect 351638 824 351644 836
rect 351696 824 351702 876
rect 368750 824 368756 876
rect 368808 864 368814 876
rect 373902 864 373908 876
rect 368808 836 373908 864
rect 368808 824 368814 836
rect 373902 824 373908 836
rect 373960 824 373966 876
rect 448238 824 448244 876
rect 448296 864 448302 876
rect 459186 864 459192 876
rect 448296 836 459192 864
rect 448296 824 448302 836
rect 459186 824 459192 836
rect 459244 824 459250 876
rect 485682 824 485688 876
rect 485740 864 485746 876
rect 498930 864 498936 876
rect 485740 836 498936 864
rect 485740 824 485746 836
rect 498930 824 498936 836
rect 498988 824 498994 876
rect 527726 824 527732 876
rect 527784 864 527790 876
rect 544378 864 544384 876
rect 527784 836 544384 864
rect 527784 824 527790 836
rect 544378 824 544384 836
rect 544436 824 544442 876
rect 547598 824 547604 876
rect 547656 864 547662 876
rect 565630 864 565636 876
rect 547656 836 565636 864
rect 547656 824 547662 836
rect 565630 824 565636 836
rect 565688 824 565694 876
rect 18230 756 18236 808
rect 18288 796 18294 808
rect 36354 796 36360 808
rect 18288 768 36360 796
rect 18288 756 18294 768
rect 36354 756 36360 768
rect 36412 756 36418 808
rect 251174 756 251180 808
rect 251232 796 251238 808
rect 253842 796 253848 808
rect 251232 768 253848 796
rect 251232 756 251238 768
rect 253842 756 253848 768
rect 253900 756 253906 808
rect 427262 756 427268 808
rect 427320 796 427326 808
rect 436738 796 436744 808
rect 427320 768 436744 796
rect 427320 756 427326 768
rect 436738 756 436744 768
rect 436796 756 436802 808
rect 442718 756 442724 808
rect 442776 796 442782 808
rect 453298 796 453304 808
rect 442776 768 453304 796
rect 442776 756 442782 768
rect 453298 756 453304 768
rect 453356 756 453362 808
rect 462406 796 462412 808
rect 460906 768 462412 796
rect 9950 688 9956 740
rect 10008 728 10014 740
rect 28626 728 28632 740
rect 10008 700 28632 728
rect 10008 688 10014 700
rect 28626 688 28632 700
rect 28684 688 28690 740
rect 401870 688 401876 740
rect 401928 728 401934 740
rect 409230 728 409236 740
rect 401928 700 409236 728
rect 401928 688 401934 700
rect 409230 688 409236 700
rect 409288 688 409294 740
rect 429470 688 429476 740
rect 429528 728 429534 740
rect 439130 728 439136 740
rect 429528 700 439136 728
rect 429528 688 429534 700
rect 439130 688 439136 700
rect 439188 688 439194 740
rect 440510 688 440516 740
rect 440568 728 440574 740
rect 450906 728 450912 740
rect 440568 700 450912 728
rect 440568 688 440574 700
rect 450906 688 450912 700
rect 450964 688 450970 740
rect 451550 688 451556 740
rect 451608 728 451614 740
rect 460906 728 460934 768
rect 462406 756 462412 768
rect 462464 756 462470 808
rect 483566 756 483572 808
rect 483624 796 483630 808
rect 497090 796 497096 808
rect 483624 768 497096 796
rect 483624 756 483630 768
rect 497090 756 497096 768
rect 497148 756 497154 808
rect 499022 756 499028 808
rect 499080 796 499086 808
rect 513558 796 513564 808
rect 499080 768 513564 796
rect 499080 756 499086 768
rect 513558 756 513564 768
rect 513616 756 513622 808
rect 528830 756 528836 808
rect 528888 796 528894 808
rect 545482 796 545488 808
rect 528888 768 545488 796
rect 528888 756 528894 768
rect 545482 756 545488 768
rect 545540 756 545546 808
rect 550910 756 550916 808
rect 550968 796 550974 808
rect 569126 796 569132 808
rect 550968 768 569132 796
rect 550968 756 550974 768
rect 569126 756 569132 768
rect 569184 756 569190 808
rect 451608 700 460934 728
rect 451608 688 451614 700
rect 468110 688 468116 740
rect 468168 728 468174 740
rect 480530 728 480536 740
rect 468168 700 480536 728
rect 468168 688 468174 700
rect 480530 688 480536 700
rect 480588 688 480594 740
rect 482462 688 482468 740
rect 482520 728 482526 740
rect 495526 728 495532 740
rect 482520 700 495532 728
rect 482520 688 482526 700
rect 495526 688 495532 700
rect 495584 688 495590 740
rect 502242 688 502248 740
rect 502300 728 502306 740
rect 517146 728 517152 740
rect 502300 700 517152 728
rect 502300 688 502306 700
rect 517146 688 517152 700
rect 517204 688 517210 740
rect 521102 688 521108 740
rect 521160 728 521166 740
rect 537202 728 537208 740
rect 521160 700 537208 728
rect 521160 688 521166 700
rect 537202 688 537208 700
rect 537260 688 537266 740
rect 537662 688 537668 740
rect 537720 728 537726 740
rect 554958 728 554964 740
rect 537720 700 554964 728
rect 537720 688 537726 700
rect 554958 688 554964 700
rect 555016 688 555022 740
rect 8754 620 8760 672
rect 8812 660 8818 672
rect 27522 660 27528 672
rect 8812 632 27528 660
rect 8812 620 8818 632
rect 27522 620 27528 632
rect 27580 620 27586 672
rect 34790 620 34796 672
rect 34848 660 34854 672
rect 51810 660 51816 672
rect 34848 632 51816 660
rect 34848 620 34854 632
rect 51810 620 51816 632
rect 51868 620 51874 672
rect 393038 620 393044 672
rect 393096 660 393102 672
rect 400122 660 400128 672
rect 393096 632 400128 660
rect 393096 620 393102 632
rect 400122 620 400128 632
rect 400180 620 400186 672
rect 400766 620 400772 672
rect 400824 660 400830 672
rect 408586 660 408592 672
rect 400824 632 408592 660
rect 400824 620 400830 632
rect 408586 620 408592 632
rect 408644 620 408650 672
rect 409598 620 409604 672
rect 409656 660 409662 672
rect 417878 660 417884 672
rect 409656 632 417884 660
rect 409656 620 409662 632
rect 417878 620 417884 632
rect 417936 620 417942 672
rect 441522 660 441528 672
rect 431926 632 441528 660
rect 14734 552 14740 604
rect 14792 552 14798 604
rect 17034 552 17040 604
rect 17092 592 17098 604
rect 35250 592 35256 604
rect 17092 564 35256 592
rect 17092 552 17098 564
rect 35250 552 35256 564
rect 35308 552 35314 604
rect 35986 552 35992 604
rect 36044 592 36050 604
rect 52914 592 52920 604
rect 36044 564 52920 592
rect 36044 552 36050 564
rect 52914 552 52920 564
rect 52972 552 52978 604
rect 389726 552 389732 604
rect 389784 592 389790 604
rect 396534 592 396540 604
rect 389784 564 396540 592
rect 389784 552 389790 564
rect 396534 552 396540 564
rect 396592 552 396598 604
rect 408402 552 408408 604
rect 408460 592 408466 604
rect 416682 592 416688 604
rect 408460 564 416688 592
rect 408460 552 408466 564
rect 416682 552 416688 564
rect 416740 552 416746 604
rect 431678 552 431684 604
rect 431736 592 431742 604
rect 431926 592 431954 632
rect 441522 620 441528 632
rect 441580 620 441586 672
rect 456978 620 456984 672
rect 457036 660 457042 672
rect 460014 660 460020 672
rect 457036 632 460020 660
rect 457036 620 457042 632
rect 460014 620 460020 632
rect 460072 620 460078 672
rect 464798 620 464804 672
rect 464856 660 464862 672
rect 476942 660 476948 672
rect 464856 632 476948 660
rect 464856 620 464862 632
rect 476942 620 476948 632
rect 477000 620 477006 672
rect 486878 620 486884 672
rect 486936 660 486942 672
rect 500586 660 500592 672
rect 486936 632 500592 660
rect 486936 620 486942 632
rect 500586 620 500592 632
rect 500644 620 500650 672
rect 503438 620 503444 672
rect 503496 660 503502 672
rect 518342 660 518348 672
rect 503496 632 518348 660
rect 503496 620 503502 632
rect 518342 620 518348 632
rect 518400 620 518406 672
rect 523310 620 523316 672
rect 523368 660 523374 672
rect 523368 632 524276 660
rect 523368 620 523374 632
rect 440326 592 440332 604
rect 431736 564 431954 592
rect 438596 564 440332 592
rect 431736 552 431742 564
rect 14752 524 14780 552
rect 33042 524 33048 536
rect 14752 496 33048 524
rect 33042 484 33048 496
rect 33100 484 33106 536
rect 39758 484 39764 536
rect 39816 524 39822 536
rect 56226 524 56232 536
rect 39816 496 56232 524
rect 39816 484 39822 496
rect 56226 484 56232 496
rect 56284 484 56290 536
rect 430482 484 430488 536
rect 430540 524 430546 536
rect 438596 524 438624 564
rect 440326 552 440332 564
rect 440384 552 440390 604
rect 447042 552 447048 604
rect 447100 592 447106 604
rect 458082 592 458088 604
rect 447100 564 458088 592
rect 447100 552 447106 564
rect 458082 552 458088 564
rect 458140 552 458146 604
rect 461486 552 461492 604
rect 461544 592 461550 604
rect 473446 592 473452 604
rect 461544 564 473452 592
rect 461544 552 461550 564
rect 473446 552 473452 564
rect 473504 552 473510 604
rect 486418 552 486424 604
rect 486476 552 486482 604
rect 498194 592 498200 604
rect 489886 564 498200 592
rect 430540 496 438624 524
rect 430540 484 430546 496
rect 459462 484 459468 536
rect 459520 524 459526 536
rect 470778 524 470784 536
rect 459520 496 470784 524
rect 459520 484 459526 496
rect 470778 484 470784 496
rect 470836 484 470842 536
rect 473630 484 473636 536
rect 473688 524 473694 536
rect 486436 524 486464 552
rect 473688 496 486464 524
rect 473688 484 473694 496
rect 16206 416 16212 468
rect 16264 456 16270 468
rect 34146 456 34152 468
rect 16264 428 34152 456
rect 16264 416 16270 428
rect 34146 416 34152 428
rect 34204 416 34210 468
rect 38562 416 38568 468
rect 38620 456 38626 468
rect 55122 456 55128 468
rect 38620 428 55128 456
rect 38620 416 38626 428
rect 55122 416 55128 428
rect 55180 416 55186 468
rect 381998 416 382004 468
rect 382056 456 382062 468
rect 387886 456 387892 468
rect 382056 428 387892 456
rect 382056 416 382062 428
rect 387886 416 387892 428
rect 387944 416 387950 468
rect 412082 416 412088 468
rect 412140 456 412146 468
rect 420362 456 420368 468
rect 412140 428 420368 456
rect 412140 416 412146 428
rect 420362 416 420368 428
rect 420420 416 420426 468
rect 437198 416 437204 468
rect 437256 456 437262 468
rect 447226 456 447232 468
rect 437256 428 447232 456
rect 437256 416 437262 428
rect 447226 416 447232 428
rect 447284 416 447290 468
rect 470318 416 470324 468
rect 470376 456 470382 468
rect 482462 456 482468 468
rect 470376 428 482468 456
rect 470376 416 470382 428
rect 482462 416 482468 428
rect 482520 416 482526 468
rect 484670 416 484676 468
rect 484728 456 484734 468
rect 489886 456 489914 564
rect 498194 552 498200 564
rect 498252 552 498258 604
rect 503806 592 503812 604
rect 498396 564 503812 592
rect 484728 428 489914 456
rect 484728 416 484734 428
rect 490190 416 490196 468
rect 490248 456 490254 468
rect 498396 456 498424 564
rect 503806 552 503812 564
rect 503864 552 503870 604
rect 508958 552 508964 604
rect 509016 592 509022 604
rect 523862 592 523868 604
rect 509016 564 523868 592
rect 509016 552 509022 564
rect 523862 552 523868 564
rect 523920 552 523926 604
rect 524248 592 524276 632
rect 524322 620 524328 672
rect 524380 660 524386 672
rect 533246 660 533252 672
rect 524380 632 533252 660
rect 524380 620 524386 632
rect 533246 620 533252 632
rect 533304 620 533310 672
rect 539594 660 539600 672
rect 533356 632 539600 660
rect 533356 592 533384 632
rect 539594 620 539600 632
rect 539652 620 539658 672
rect 542078 620 542084 672
rect 542136 660 542142 672
rect 542136 632 544976 660
rect 542136 620 542142 632
rect 524248 564 533384 592
rect 533706 552 533712 604
rect 533764 552 533770 604
rect 533798 552 533804 604
rect 533856 592 533862 604
rect 533856 564 543044 592
rect 533856 552 533862 564
rect 512086 524 512092 536
rect 490248 428 498424 456
rect 499546 496 512092 524
rect 490248 416 490254 428
rect 11514 348 11520 400
rect 11572 388 11578 400
rect 29730 388 29736 400
rect 11572 360 29736 388
rect 11572 348 11578 360
rect 29730 348 29736 360
rect 29788 348 29794 400
rect 32214 348 32220 400
rect 32272 388 32278 400
rect 49602 388 49608 400
rect 32272 360 49608 388
rect 32272 348 32278 360
rect 49602 348 49608 360
rect 49660 348 49666 400
rect 407390 348 407396 400
rect 407448 388 407454 400
rect 415302 388 415308 400
rect 407448 360 415308 388
rect 407448 348 407454 360
rect 415302 348 415308 360
rect 415360 348 415366 400
rect 460566 348 460572 400
rect 460624 388 460630 400
rect 472434 388 472440 400
rect 460624 360 472440 388
rect 460624 348 460630 360
rect 472434 348 472440 360
rect 472492 348 472498 400
rect 478322 348 478328 400
rect 478380 388 478386 400
rect 490742 388 490748 400
rect 478380 360 490748 388
rect 478380 348 478386 360
rect 490742 348 490748 360
rect 490800 348 490806 400
rect 497918 348 497924 400
rect 497976 388 497982 400
rect 499546 388 499574 496
rect 512086 484 512092 496
rect 512144 484 512150 536
rect 517790 484 517796 536
rect 517848 524 517854 536
rect 533724 524 533752 552
rect 517848 496 533752 524
rect 517848 484 517854 496
rect 500126 416 500132 468
rect 500184 456 500190 468
rect 514938 456 514944 468
rect 500184 428 514944 456
rect 500184 416 500190 428
rect 514938 416 514944 428
rect 514996 416 515002 468
rect 525702 416 525708 468
rect 525760 456 525766 468
rect 542170 456 542176 468
rect 525760 428 542176 456
rect 525760 416 525766 428
rect 542170 416 542176 428
rect 542228 416 542234 468
rect 497976 360 499574 388
rect 497976 348 497982 360
rect 504542 348 504548 400
rect 504600 388 504606 400
rect 519722 388 519728 400
rect 504600 360 519728 388
rect 504600 348 504606 360
rect 519722 348 519728 360
rect 519780 348 519786 400
rect 533246 348 533252 400
rect 533304 388 533310 400
rect 540422 388 540428 400
rect 533304 360 540428 388
rect 533304 348 533310 360
rect 540422 348 540428 360
rect 540480 348 540486 400
rect 543016 388 543044 564
rect 544948 524 544976 632
rect 548978 620 548984 672
rect 549036 660 549042 672
rect 566826 660 566832 672
rect 549036 632 566832 660
rect 549036 620 549042 632
rect 566826 620 566832 632
rect 566884 620 566890 672
rect 545390 552 545396 604
rect 545448 592 545454 604
rect 563238 592 563244 604
rect 545448 564 563244 592
rect 545448 552 545454 564
rect 563238 552 563244 564
rect 563296 552 563302 604
rect 559374 524 559380 536
rect 544948 496 559380 524
rect 559374 484 559380 496
rect 559432 484 559438 536
rect 544562 416 544568 468
rect 544620 456 544626 468
rect 562226 456 562232 468
rect 544620 428 562232 456
rect 544620 416 544626 428
rect 562226 416 562232 428
rect 562284 416 562290 468
rect 550450 388 550456 400
rect 543016 360 550456 388
rect 550450 348 550456 360
rect 550508 348 550514 400
rect 555326 348 555332 400
rect 555384 388 555390 400
rect 573542 388 573548 400
rect 555384 360 573548 388
rect 555384 348 555390 360
rect 573542 348 573548 360
rect 573600 348 573606 400
rect 3234 280 3240 332
rect 3292 320 3298 332
rect 22002 320 22008 332
rect 3292 292 22008 320
rect 3292 280 3298 292
rect 22002 280 22008 292
rect 22060 280 22066 332
rect 30282 280 30288 332
rect 30340 320 30346 332
rect 47394 320 47400 332
rect 30340 292 47400 320
rect 30340 280 30346 292
rect 47394 280 47400 292
rect 47452 280 47458 332
rect 398558 280 398564 332
rect 398616 320 398622 332
rect 406194 320 406200 332
rect 398616 292 406200 320
rect 398616 280 398622 292
rect 406194 280 406200 292
rect 406252 280 406258 332
rect 410978 280 410984 332
rect 411036 320 411042 332
rect 418614 320 418620 332
rect 411036 292 418620 320
rect 411036 280 411042 292
rect 418614 280 418620 292
rect 418672 280 418678 332
rect 453758 280 453764 332
rect 453816 320 453822 332
rect 464982 320 464988 332
rect 453816 292 464988 320
rect 453816 280 453822 292
rect 464982 280 464988 292
rect 465040 280 465046 332
rect 471422 280 471428 332
rect 471480 320 471486 332
rect 484210 320 484216 332
rect 471480 292 484216 320
rect 471480 280 471486 292
rect 484210 280 484216 292
rect 484268 280 484274 332
rect 505646 280 505652 332
rect 505704 320 505710 332
rect 520366 320 520372 332
rect 505704 292 520372 320
rect 505704 280 505710 292
rect 520366 280 520372 292
rect 520424 280 520430 332
rect 531038 280 531044 332
rect 531096 320 531102 332
rect 548058 320 548064 332
rect 531096 292 548064 320
rect 531096 280 531102 292
rect 548058 280 548064 292
rect 548116 280 548122 332
rect 551922 280 551928 332
rect 551980 320 551986 332
rect 570506 320 570512 332
rect 551980 292 570512 320
rect 551980 280 551986 292
rect 570506 280 570512 292
rect 570564 280 570570 332
rect 22830 212 22836 264
rect 22888 252 22894 264
rect 40494 252 40500 264
rect 22888 224 40500 252
rect 22888 212 22894 224
rect 40494 212 40500 224
rect 40552 212 40558 264
rect 42242 212 42248 264
rect 42300 252 42306 264
rect 58158 252 58164 264
rect 42300 224 58164 252
rect 42300 212 42306 224
rect 58158 212 58164 224
rect 58216 212 58222 264
rect 354398 212 354404 264
rect 354456 252 354462 264
rect 358906 252 358912 264
rect 354456 224 358912 252
rect 354456 212 354462 224
rect 358906 212 358912 224
rect 358964 212 358970 264
rect 380802 212 380808 264
rect 380860 252 380866 264
rect 386782 252 386788 264
rect 380860 224 386788 252
rect 380860 212 380866 224
rect 386782 212 386788 224
rect 386840 212 386846 264
rect 391658 212 391664 264
rect 391716 252 391722 264
rect 398742 252 398748 264
rect 391716 224 398748 252
rect 391716 212 391722 224
rect 398742 212 398748 224
rect 398800 212 398806 264
rect 405182 212 405188 264
rect 405240 252 405246 264
rect 412818 252 412824 264
rect 405240 224 412824 252
rect 405240 212 405246 224
rect 412818 212 412824 224
rect 412876 212 412882 264
rect 457898 212 457904 264
rect 457956 252 457962 264
rect 470042 252 470048 264
rect 457956 224 470048 252
rect 457956 212 457962 224
rect 470042 212 470048 224
rect 470100 212 470106 264
rect 472526 212 472532 264
rect 472584 252 472590 264
rect 484854 252 484860 264
rect 472584 224 484860 252
rect 472584 212 472590 224
rect 484854 212 484860 224
rect 484912 212 484918 264
rect 511442 212 511448 264
rect 511500 252 511506 264
rect 526254 252 526260 264
rect 511500 224 526260 252
rect 511500 212 511506 224
rect 526254 212 526260 224
rect 526312 212 526318 264
rect 538766 212 538772 264
rect 538824 252 538830 264
rect 556338 252 556344 264
rect 538824 224 556344 252
rect 538824 212 538830 224
rect 556338 212 556344 224
rect 556396 212 556402 264
rect 557166 212 557172 264
rect 557224 252 557230 264
rect 575934 252 575940 264
rect 557224 224 575940 252
rect 557224 212 557230 224
rect 575934 212 575940 224
rect 575992 212 575998 264
rect 8018 144 8024 196
rect 8076 184 8082 196
rect 26326 184 26332 196
rect 8076 156 26332 184
rect 8076 144 8082 156
rect 26326 144 26332 156
rect 26384 144 26390 196
rect 31110 144 31116 196
rect 31168 184 31174 196
rect 48498 184 48504 196
rect 31168 156 48504 184
rect 31168 144 31174 156
rect 48498 144 48504 156
rect 48556 144 48562 196
rect 53558 144 53564 196
rect 53616 184 53622 196
rect 69474 184 69480 196
rect 53616 156 69480 184
rect 53616 144 53622 156
rect 69474 144 69480 156
rect 69532 144 69538 196
rect 418430 144 418436 196
rect 418488 184 418494 196
rect 426894 184 426900 196
rect 418488 156 426900 184
rect 418488 144 418494 156
rect 426894 144 426900 156
rect 426952 144 426958 196
rect 465810 144 465816 196
rect 465868 184 465874 196
rect 478322 184 478328 196
rect 465868 156 478328 184
rect 465868 144 465874 156
rect 478322 144 478328 156
rect 478380 144 478386 196
rect 479150 144 479156 196
rect 479208 184 479214 196
rect 492490 184 492496 196
rect 479208 156 492496 184
rect 479208 144 479214 156
rect 492490 144 492496 156
rect 492548 144 492554 196
rect 492582 144 492588 196
rect 492640 184 492646 196
rect 506658 184 506664 196
rect 492640 156 506664 184
rect 492640 144 492646 156
rect 506658 144 506664 156
rect 506716 144 506722 196
rect 512638 144 512644 196
rect 512696 184 512702 196
rect 528002 184 528008 196
rect 512696 156 528008 184
rect 512696 144 512702 156
rect 528002 144 528008 156
rect 528060 144 528066 196
rect 535362 144 535368 196
rect 535420 184 535426 196
rect 552842 184 552848 196
rect 535420 156 552848 184
rect 535420 144 535426 156
rect 552842 144 552848 156
rect 552900 144 552906 196
rect 554222 144 554228 196
rect 554280 184 554286 196
rect 572898 184 572904 196
rect 554280 156 572904 184
rect 554280 144 554286 156
rect 572898 144 572904 156
rect 572956 144 572962 196
rect 22002 76 22008 128
rect 22060 116 22066 128
rect 39390 116 39396 128
rect 22060 88 39396 116
rect 22060 76 22066 88
rect 39390 76 39396 88
rect 39448 76 39454 128
rect 45278 76 45284 128
rect 45336 116 45342 128
rect 61746 116 61752 128
rect 45336 88 61752 116
rect 45336 76 45342 88
rect 61746 76 61752 88
rect 61804 76 61810 128
rect 399662 76 399668 128
rect 399720 116 399726 128
rect 407022 116 407028 128
rect 399720 88 407028 116
rect 399720 76 399726 88
rect 407022 76 407028 88
rect 407080 76 407086 128
rect 423950 76 423956 128
rect 424008 116 424014 128
rect 433426 116 433432 128
rect 424008 88 433432 116
rect 424008 76 424014 88
rect 433426 76 433432 88
rect 433484 76 433490 128
rect 452562 76 452568 128
rect 452620 116 452626 128
rect 464154 116 464160 128
rect 452620 88 464160 116
rect 452620 76 452626 88
rect 464154 76 464160 88
rect 464212 76 464218 128
rect 467006 76 467012 128
rect 467064 116 467070 128
rect 478966 116 478972 128
rect 467064 88 478972 116
rect 467064 76 467070 88
rect 478966 76 478972 88
rect 479024 76 479030 128
rect 491294 76 491300 128
rect 491352 116 491358 128
rect 505554 116 505560 128
rect 491352 88 505560 116
rect 491352 76 491358 88
rect 505554 76 505560 88
rect 505612 76 505618 128
rect 514478 76 514484 128
rect 514536 116 514542 128
rect 529934 116 529940 128
rect 514536 88 529940 116
rect 514536 76 514542 88
rect 529934 76 529940 88
rect 529992 76 529998 128
rect 540974 76 540980 128
rect 541032 116 541038 128
rect 558730 116 558736 128
rect 541032 88 558736 116
rect 541032 76 541038 88
rect 558730 76 558736 88
rect 558788 76 558794 128
rect 558822 76 558828 128
rect 558880 116 558886 128
rect 577130 116 577136 128
rect 558880 88 577136 116
rect 558880 76 558886 88
rect 577130 76 577136 88
rect 577188 76 577194 128
rect 382 8 388 60
rect 440 48 446 60
rect 19794 48 19800 60
rect 440 20 19800 48
rect 440 8 446 20
rect 19794 8 19800 20
rect 19852 8 19858 60
rect 24578 8 24584 60
rect 24636 48 24642 60
rect 41598 48 41604 60
rect 24636 20 41604 48
rect 24636 8 24642 20
rect 41598 8 41604 20
rect 41656 8 41662 60
rect 42886 8 42892 60
rect 42944 48 42950 60
rect 59354 48 59360 60
rect 42944 20 59360 48
rect 42944 8 42950 20
rect 59354 8 59360 20
rect 59412 8 59418 60
rect 344738 8 344744 60
rect 344796 48 344802 60
rect 348234 48 348240 60
rect 344796 20 348240 48
rect 344796 8 344802 20
rect 348234 8 348240 20
rect 348292 8 348298 60
rect 363230 8 363236 60
rect 363288 48 363294 60
rect 367830 48 367836 60
rect 363288 20 367836 48
rect 363288 8 363294 20
rect 367830 8 367836 20
rect 367888 8 367894 60
rect 383102 8 383108 60
rect 383160 48 383166 60
rect 389634 48 389640 60
rect 383160 20 389640 48
rect 383160 8 383166 20
rect 389634 8 389640 20
rect 389692 8 389698 60
rect 390830 8 390836 60
rect 390888 48 390894 60
rect 397914 48 397920 60
rect 390888 20 397920 48
rect 390888 8 390894 20
rect 397914 8 397920 20
rect 397972 8 397978 60
rect 402882 8 402888 60
rect 402940 48 402946 60
rect 410978 48 410984 60
rect 402940 20 410984 48
rect 402940 8 402946 20
rect 410978 8 410984 20
rect 411036 8 411042 60
rect 417326 8 417332 60
rect 417384 48 417390 60
rect 425790 48 425796 60
rect 417384 20 425796 48
rect 417384 8 417390 20
rect 425790 8 425796 20
rect 425848 8 425854 60
rect 463602 8 463608 60
rect 463660 48 463666 60
rect 475930 48 475936 60
rect 463660 20 475936 48
rect 463660 8 463666 20
rect 475930 8 475936 20
rect 475988 8 475994 60
rect 477218 8 477224 60
rect 477276 48 477282 60
rect 490098 48 490104 60
rect 477276 20 490104 48
rect 477276 8 477282 20
rect 490098 8 490104 20
rect 490156 8 490162 60
rect 496722 8 496728 60
rect 496780 48 496786 60
rect 511442 48 511448 60
rect 496780 20 511448 48
rect 496780 8 496786 20
rect 511442 8 511448 20
rect 511500 8 511506 60
rect 526898 8 526904 60
rect 526956 48 526962 60
rect 542814 48 542820 60
rect 526956 20 542820 48
rect 526956 8 526962 20
rect 542814 8 542820 20
rect 542872 8 542878 60
rect 546402 8 546408 60
rect 546460 48 546466 60
rect 564618 48 564624 60
rect 546460 20 564624 48
rect 546460 8 546466 20
rect 564618 8 564624 20
rect 564676 8 564682 60
<< via1 >>
rect 186504 702992 186556 703044
rect 188436 702992 188488 703044
rect 235172 702992 235224 703044
rect 236184 702992 236236 703044
rect 522764 702992 522816 703044
rect 527088 702992 527140 703044
rect 570512 702992 570564 703044
rect 575848 702992 575900 703044
rect 490932 702720 490984 702772
rect 494796 702720 494848 702772
rect 538680 702720 538732 702772
rect 543464 702720 543516 702772
rect 24308 702448 24360 702500
rect 29276 702448 29328 702500
rect 218980 702448 219032 702500
rect 220268 702448 220320 702500
rect 459100 702448 459152 702500
rect 462320 702448 462372 702500
rect 506848 702448 506900 702500
rect 510988 702448 511040 702500
rect 554596 702448 554648 702500
rect 559656 702448 559708 702500
rect 8116 700952 8168 701004
rect 13084 700952 13136 701004
rect 40500 700952 40552 701004
rect 44916 700952 44968 701004
rect 56784 700952 56836 701004
rect 60740 700952 60792 701004
rect 72976 700952 73028 701004
rect 76748 700952 76800 701004
rect 89168 700952 89220 701004
rect 92572 700952 92624 701004
rect 105452 700952 105504 701004
rect 108580 700952 108632 701004
rect 121644 700952 121696 701004
rect 124404 700952 124456 701004
rect 137836 700952 137888 701004
rect 140412 700952 140464 701004
rect 154120 700952 154172 701004
rect 156236 700952 156288 701004
rect 170312 700952 170364 701004
rect 172428 700952 172480 701004
rect 202788 700952 202840 701004
rect 204260 700952 204312 701004
rect 348056 700952 348108 701004
rect 348792 700952 348844 701004
rect 363880 700952 363932 701004
rect 364984 700952 365036 701004
rect 379336 700952 379388 701004
rect 381176 700952 381228 701004
rect 395712 700952 395764 701004
rect 397460 700952 397512 701004
rect 411720 700952 411772 701004
rect 413652 700952 413704 701004
rect 427544 700952 427596 701004
rect 429844 700952 429896 701004
rect 443552 700952 443604 701004
rect 446128 700952 446180 701004
rect 475384 700952 475436 701004
rect 478512 700952 478564 701004
rect 59728 3816 59780 3868
rect 74724 3952 74776 4004
rect 58808 3680 58860 3732
rect 70216 3884 70268 3936
rect 62028 3748 62080 3800
rect 67456 3748 67508 3800
rect 78036 3884 78088 3936
rect 63224 3612 63276 3664
rect 69020 3680 69072 3732
rect 71412 3680 71464 3732
rect 69112 3612 69164 3664
rect 83556 3816 83608 3868
rect 80888 3748 80940 3800
rect 94596 3816 94648 3868
rect 122288 3816 122340 3868
rect 133236 3816 133288 3868
rect 84476 3748 84528 3800
rect 98000 3748 98052 3800
rect 114008 3748 114060 3800
rect 125508 3748 125560 3800
rect 66720 3544 66772 3596
rect 81348 3680 81400 3732
rect 85672 3680 85724 3732
rect 56048 3476 56100 3528
rect 69020 3476 69072 3528
rect 70124 3476 70176 3528
rect 54944 3408 54996 3460
rect 70216 3408 70268 3460
rect 72976 3476 73028 3528
rect 86868 3612 86920 3664
rect 87788 3680 87840 3732
rect 101220 3680 101272 3732
rect 116400 3680 116452 3732
rect 127716 3680 127768 3732
rect 99012 3612 99064 3664
rect 109408 3612 109460 3664
rect 121184 3612 121236 3664
rect 125048 3612 125100 3664
rect 135444 3612 135496 3664
rect 143632 3612 143684 3664
rect 153108 3612 153160 3664
rect 82912 3544 82964 3596
rect 83280 3544 83332 3596
rect 96804 3544 96856 3596
rect 102232 3544 102284 3596
rect 114468 3544 114520 3596
rect 121092 3544 121144 3596
rect 132132 3544 132184 3596
rect 136456 3544 136508 3596
rect 146484 3544 146536 3596
rect 149520 3544 149572 3596
rect 158628 3544 158680 3596
rect 78588 3476 78640 3528
rect 92388 3476 92440 3528
rect 51356 3340 51408 3392
rect 66996 3340 67048 3392
rect 67456 3340 67508 3392
rect 76932 3340 76984 3392
rect 65524 3272 65576 3324
rect 50160 3204 50212 3256
rect 65892 3204 65944 3256
rect 71504 3272 71556 3324
rect 85764 3408 85816 3460
rect 90364 3408 90416 3460
rect 103612 3476 103664 3528
rect 110512 3476 110564 3528
rect 122380 3476 122432 3528
rect 127072 3476 127124 3528
rect 137652 3476 137704 3528
rect 139216 3476 139268 3528
rect 148692 3476 148744 3528
rect 153016 3476 153068 3528
rect 160192 3476 160244 3528
rect 79692 3340 79744 3392
rect 83004 3340 83056 3392
rect 89536 3340 89588 3392
rect 102324 3408 102376 3460
rect 105728 3408 105780 3460
rect 117780 3408 117832 3460
rect 131764 3408 131816 3460
rect 142252 3408 142304 3460
rect 142528 3408 142580 3460
rect 151728 3408 151780 3460
rect 155776 3408 155828 3460
rect 96252 3340 96304 3392
rect 109040 3340 109092 3392
rect 112812 3340 112864 3392
rect 124128 3340 124180 3392
rect 125968 3340 126020 3392
rect 136640 3340 136692 3392
rect 82912 3272 82964 3324
rect 84660 3272 84712 3324
rect 86868 3272 86920 3324
rect 100116 3272 100168 3324
rect 103336 3272 103388 3324
rect 115572 3272 115624 3324
rect 117596 3272 117648 3324
rect 128820 3272 128872 3324
rect 129372 3272 129424 3324
rect 139860 3272 139912 3324
rect 149796 3340 149848 3392
rect 148324 3272 148376 3324
rect 157248 3272 157300 3324
rect 79968 3204 80020 3256
rect 93952 3204 94004 3256
rect 106740 3204 106792 3256
rect 107200 3204 107252 3256
rect 118608 3204 118660 3256
rect 119896 3204 119948 3256
rect 131028 3204 131080 3256
rect 140044 3204 140096 3256
rect 154028 3204 154080 3256
rect 40960 3136 41012 3188
rect 57060 3136 57112 3188
rect 57520 3136 57572 3188
rect 72516 3136 72568 3188
rect 73804 3136 73856 3188
rect 87972 3136 88024 3188
rect 101036 3136 101088 3188
rect 113088 3136 113140 3188
rect 52552 3068 52604 3120
rect 68100 3068 68152 3120
rect 76288 3068 76340 3120
rect 44272 3000 44324 3052
rect 60372 3000 60424 3052
rect 64328 3000 64380 3052
rect 79140 3000 79192 3052
rect 79600 3068 79652 3120
rect 89076 3068 89128 3120
rect 98736 3068 98788 3120
rect 111156 3068 111208 3120
rect 111616 3068 111668 3120
rect 123300 3068 123352 3120
rect 33600 2932 33652 2984
rect 50436 2932 50488 2984
rect 26608 2864 26660 2916
rect 43812 2864 43864 2916
rect 48964 2864 49016 2916
rect 64880 2932 64932 2984
rect 67916 2932 67968 2984
rect 82728 2932 82780 2984
rect 83004 3000 83056 3052
rect 93492 3000 93544 3052
rect 95148 3000 95200 3052
rect 107844 3000 107896 3052
rect 108488 3000 108540 3052
rect 119988 3000 120040 3052
rect 134340 3136 134392 3188
rect 137652 3136 137704 3188
rect 147772 3136 147824 3188
rect 134156 3068 134208 3120
rect 144276 3068 144328 3120
rect 147128 3068 147180 3120
rect 156420 3136 156472 3188
rect 128176 3000 128228 3052
rect 138756 3000 138808 3052
rect 90456 2932 90508 2984
rect 91560 2932 91612 2984
rect 104532 2932 104584 2984
rect 104624 2932 104676 2984
rect 116952 2932 117004 2984
rect 123484 2932 123536 2984
rect 130568 2932 130620 2984
rect 140964 2932 141016 2984
rect 27712 2796 27764 2848
rect 45192 2796 45244 2848
rect 47860 2796 47912 2848
rect 63684 2864 63736 2916
rect 75368 2864 75420 2916
rect 79600 2864 79652 2916
rect 82084 2864 82136 2916
rect 95976 2864 96028 2916
rect 97448 2864 97500 2916
rect 110052 2864 110104 2916
rect 115204 2864 115256 2916
rect 126888 2864 126940 2916
rect 132960 2864 133012 2916
rect 143172 3000 143224 3052
rect 145932 3000 145984 3052
rect 155316 3068 155368 3120
rect 166080 3408 166132 3460
rect 158168 3272 158220 3324
rect 166356 3340 166408 3392
rect 174084 3340 174136 3392
rect 161296 3272 161348 3324
rect 169668 3272 169720 3324
rect 181812 3272 181864 3324
rect 564348 3272 564400 3324
rect 583392 3272 583444 3324
rect 160192 3204 160244 3256
rect 161940 3204 161992 3256
rect 163688 3204 163740 3256
rect 171876 3204 171928 3256
rect 174268 3204 174320 3256
rect 164148 3136 164200 3188
rect 170772 3136 170824 3188
rect 178500 3136 178552 3188
rect 162768 3068 162820 3120
rect 164884 3068 164936 3120
rect 172980 3068 173032 3120
rect 173440 3068 173492 3120
rect 180892 3204 180944 3256
rect 184940 3204 184992 3256
rect 181444 3136 181496 3188
rect 188436 3136 188488 3188
rect 200304 3204 200356 3256
rect 206100 3204 206152 3256
rect 556712 3204 556764 3256
rect 575112 3204 575164 3256
rect 191748 3136 191800 3188
rect 195612 3136 195664 3188
rect 201684 3136 201736 3188
rect 220268 3136 220320 3188
rect 224868 3136 224920 3188
rect 561128 3136 561180 3188
rect 579804 3136 579856 3188
rect 179052 3068 179104 3120
rect 186320 3068 186372 3120
rect 190552 3068 190604 3120
rect 197268 3068 197320 3120
rect 202696 3068 202748 3120
rect 208308 3068 208360 3120
rect 209872 3068 209924 3120
rect 214932 3068 214984 3120
rect 215668 3068 215720 3120
rect 220452 3068 220504 3120
rect 221556 3068 221608 3120
rect 225972 3068 226024 3120
rect 228732 3068 228784 3120
rect 232596 3068 232648 3120
rect 239312 3068 239364 3120
rect 242532 3068 242584 3120
rect 543464 3068 543516 3120
rect 560484 3068 560536 3120
rect 562232 3068 562284 3120
rect 581000 3068 581052 3120
rect 151820 3000 151872 3052
rect 160836 3000 160888 3052
rect 162492 3000 162544 3052
rect 170864 3000 170916 3052
rect 171968 3000 172020 3052
rect 179604 3000 179656 3052
rect 182548 3000 182600 3052
rect 189540 3000 189592 3052
rect 189724 3000 189776 3052
rect 196164 3000 196216 3052
rect 141240 2932 141292 2984
rect 150900 2932 150952 2984
rect 156604 2932 156656 2984
rect 165528 2932 165580 2984
rect 167184 2932 167236 2984
rect 175464 2932 175516 2984
rect 175832 2932 175884 2984
rect 144736 2864 144788 2916
rect 60832 2796 60884 2848
rect 75828 2796 75880 2848
rect 77392 2796 77444 2848
rect 91284 2796 91336 2848
rect 92756 2796 92808 2848
rect 98644 2796 98696 2848
rect 99840 2796 99892 2848
rect 112536 2796 112588 2848
rect 118792 2796 118844 2848
rect 130200 2796 130252 2848
rect 135260 2796 135312 2848
rect 145380 2796 145432 2848
rect 150624 2864 150676 2916
rect 160008 2864 160060 2916
rect 160100 2864 160152 2916
rect 168840 2864 168892 2916
rect 169576 2864 169628 2916
rect 177672 2864 177724 2916
rect 177856 2932 177908 2984
rect 185400 2932 185452 2984
rect 194416 2932 194468 2984
rect 200580 3000 200632 3052
rect 203892 3000 203944 3052
rect 209412 3000 209464 3052
rect 212172 3000 212224 3052
rect 217140 3000 217192 3052
rect 219256 3000 219308 3052
rect 223488 3000 223540 3052
rect 228180 3000 228232 3052
rect 229836 3000 229888 3052
rect 233700 3000 233752 3052
rect 234620 3000 234672 3052
rect 238116 3000 238168 3052
rect 240508 3000 240560 3052
rect 243636 3000 243688 3052
rect 245200 3000 245252 3052
rect 248052 3000 248104 3052
rect 248788 3000 248840 3052
rect 251364 3000 251416 3052
rect 333704 3000 333756 3052
rect 336280 3000 336332 3052
rect 530032 3000 530084 3052
rect 546684 3000 546736 3052
rect 553308 3000 553360 3052
rect 571524 3000 571576 3052
rect 199108 2932 199160 2984
rect 204996 2932 205048 2984
rect 182916 2864 182968 2916
rect 183744 2864 183796 2916
rect 190644 2864 190696 2916
rect 192392 2864 192444 2916
rect 198372 2864 198424 2916
rect 201500 2864 201552 2916
rect 206928 2932 206980 2984
rect 208584 2932 208636 2984
rect 213828 2932 213880 2984
rect 214472 2932 214524 2984
rect 219348 2932 219400 2984
rect 223948 2932 224000 2984
rect 225144 2932 225196 2984
rect 229560 2932 229612 2984
rect 231032 2932 231084 2984
rect 235080 2932 235132 2984
rect 235816 2932 235868 2984
rect 239496 2932 239548 2984
rect 242072 2932 242124 2984
rect 245016 2932 245068 2984
rect 247592 2932 247644 2984
rect 250536 2932 250588 2984
rect 253480 2932 253532 2984
rect 256056 2932 256108 2984
rect 310244 2932 310296 2984
rect 311440 2932 311492 2984
rect 325700 2932 325752 2984
rect 328000 2932 328052 2984
rect 329012 2932 329064 2984
rect 331588 2932 331640 2984
rect 332324 2932 332376 2984
rect 335084 2932 335136 2984
rect 341156 2932 341208 2984
rect 344560 2932 344612 2984
rect 513288 2932 513340 2984
rect 529020 2932 529072 2984
rect 549812 2932 549864 2984
rect 568028 2932 568080 2984
rect 206192 2864 206244 2916
rect 211620 2864 211672 2916
rect 213368 2864 213420 2916
rect 217968 2864 218020 2916
rect 218060 2864 218112 2916
rect 222936 2864 222988 2916
rect 223120 2864 223172 2916
rect 227352 2864 227404 2916
rect 227536 2864 227588 2916
rect 231768 2864 231820 2916
rect 232228 2864 232280 2916
rect 236184 2864 236236 2916
rect 237012 2864 237064 2916
rect 240600 2864 240652 2916
rect 244096 2864 244148 2916
rect 247224 2864 247276 2916
rect 249984 2864 250036 2916
rect 252744 2864 252796 2916
rect 254676 2864 254728 2916
rect 257160 2864 257212 2916
rect 261760 2864 261812 2916
rect 263784 2864 263836 2916
rect 312452 2864 312504 2916
rect 313832 2864 313884 2916
rect 314568 2864 314620 2916
rect 316224 2864 316276 2916
rect 316868 2864 316920 2916
rect 318524 2864 318576 2916
rect 319076 2864 319128 2916
rect 320916 2864 320968 2916
rect 321284 2864 321336 2916
rect 323308 2864 323360 2916
rect 323492 2864 323544 2916
rect 325608 2864 325660 2916
rect 327908 2864 327960 2916
rect 330392 2864 330444 2916
rect 331128 2864 331180 2916
rect 333888 2864 333940 2916
rect 334532 2864 334584 2916
rect 337476 2864 337528 2916
rect 340052 2864 340104 2916
rect 342996 2864 343048 2916
rect 517520 2864 517572 2916
rect 523040 2864 523092 2916
rect 525800 2864 525852 2916
rect 531320 2864 531372 2916
rect 536564 2864 536616 2916
rect 553768 2864 553820 2916
rect 559748 2864 559800 2916
rect 578608 2864 578660 2916
rect 154212 2796 154264 2848
rect 158904 2796 158956 2848
rect 167736 2796 167788 2848
rect 168380 2796 168432 2848
rect 176292 2796 176344 2848
rect 180248 2796 180300 2848
rect 187332 2796 187384 2848
rect 199476 2796 199528 2848
rect 205088 2796 205140 2848
rect 210516 2796 210568 2848
rect 210976 2796 211028 2848
rect 216036 2796 216088 2848
rect 216864 2796 216916 2848
rect 221832 2796 221884 2848
rect 226340 2796 226392 2848
rect 230664 2796 230716 2848
rect 233424 2796 233476 2848
rect 237288 2796 237340 2848
rect 238116 2796 238168 2848
rect 241704 2796 241756 2848
rect 242900 2796 242952 2848
rect 246120 2796 246172 2848
rect 246396 2796 246448 2848
rect 249432 2796 249484 2848
rect 252376 2796 252428 2848
rect 254952 2796 255004 2848
rect 255872 2796 255924 2848
rect 258264 2796 258316 2848
rect 260656 2796 260708 2848
rect 262680 2796 262732 2848
rect 304724 2796 304776 2848
rect 305552 2796 305604 2848
rect 306932 2796 306984 2848
rect 307944 2796 307996 2848
rect 309140 2796 309192 2848
rect 310244 2796 310296 2848
rect 311348 2796 311400 2848
rect 312636 2796 312688 2848
rect 313556 2796 313608 2848
rect 315028 2796 315080 2848
rect 315764 2796 315816 2848
rect 317328 2796 317380 2848
rect 317972 2796 318024 2848
rect 319720 2796 319772 2848
rect 320088 2796 320140 2848
rect 322112 2796 322164 2848
rect 322388 2796 322440 2848
rect 324412 2796 324464 2848
rect 324596 2796 324648 2848
rect 326804 2796 326856 2848
rect 326988 2796 327040 2848
rect 329196 2796 329248 2848
rect 330116 2796 330168 2848
rect 332692 2796 332744 2848
rect 335636 2796 335688 2848
rect 338672 2796 338724 2848
rect 338948 2796 339000 2848
rect 342076 2796 342128 2848
rect 346676 2796 346728 2848
rect 350448 2796 350500 2848
rect 353208 2796 353260 2848
rect 357532 2796 357584 2848
rect 372344 2796 372396 2848
rect 377680 2796 377732 2848
rect 517612 2796 517664 2848
rect 521844 2796 521896 2848
rect 562968 2796 563020 2848
rect 582196 2796 582248 2848
rect 193220 2728 193272 2780
rect 176660 1300 176712 1352
rect 184296 1300 184348 1352
rect 187332 1300 187384 1352
rect 194232 1300 194284 1352
rect 198280 1300 198332 1352
rect 204168 1300 204220 1352
rect 207388 1300 207440 1352
rect 213000 1300 213052 1352
rect 257068 1300 257120 1352
rect 259368 1300 259420 1352
rect 259460 1300 259512 1352
rect 261576 1300 261628 1352
rect 262956 1300 263008 1352
rect 264888 1300 264940 1352
rect 265348 1300 265400 1352
rect 267096 1300 267148 1352
rect 267740 1300 267792 1352
rect 269304 1300 269356 1352
rect 271236 1300 271288 1352
rect 272616 1300 272668 1352
rect 273628 1300 273680 1352
rect 274824 1300 274876 1352
rect 277124 1300 277176 1352
rect 278136 1300 278188 1352
rect 279516 1300 279568 1352
rect 280344 1300 280396 1352
rect 336648 1300 336700 1352
rect 339868 1300 339920 1352
rect 342168 1300 342220 1352
rect 345756 1300 345808 1352
rect 348884 1300 348936 1352
rect 352840 1300 352892 1352
rect 356612 1300 356664 1352
rect 361120 1300 361172 1352
rect 364248 1300 364300 1352
rect 369400 1300 369452 1352
rect 374276 1300 374328 1352
rect 379612 1300 379664 1352
rect 384212 1300 384264 1352
rect 390652 1300 390704 1352
rect 396356 1300 396408 1352
rect 403624 1300 403676 1352
rect 406292 1300 406344 1352
rect 414296 1300 414348 1352
rect 419448 1300 419500 1352
rect 428280 1300 428332 1352
rect 428372 1300 428424 1352
rect 98644 1232 98696 1284
rect 105912 1232 105964 1284
rect 188896 1232 188948 1284
rect 195336 1232 195388 1284
rect 197176 1232 197228 1284
rect 203064 1232 203116 1284
rect 258264 1232 258316 1284
rect 260472 1232 260524 1284
rect 264152 1232 264204 1284
rect 265992 1232 266044 1284
rect 266544 1232 266596 1284
rect 268200 1232 268252 1284
rect 270040 1232 270092 1284
rect 271512 1232 271564 1284
rect 272432 1232 272484 1284
rect 273720 1232 273772 1284
rect 343364 1232 343416 1284
rect 346952 1232 347004 1284
rect 349988 1232 350040 1284
rect 354036 1232 354088 1284
rect 357716 1232 357768 1284
rect 362316 1232 362368 1284
rect 365444 1232 365496 1284
rect 370228 1232 370280 1284
rect 370964 1232 371016 1284
rect 376116 1232 376168 1284
rect 377588 1232 377640 1284
rect 383568 1232 383620 1284
rect 388628 1232 388680 1284
rect 395344 1232 395396 1284
rect 404084 1232 404136 1284
rect 411904 1232 411956 1284
rect 413928 1232 413980 1284
rect 422576 1232 422628 1284
rect 426164 1232 426216 1284
rect 435180 1232 435232 1284
rect 436008 1300 436060 1352
rect 437572 1232 437624 1284
rect 438308 1232 438360 1284
rect 443828 1300 443880 1352
rect 454132 1300 454184 1352
rect 186136 1164 186188 1216
rect 193128 1164 193180 1216
rect 268844 1164 268896 1216
rect 270408 1164 270460 1216
rect 359924 1164 359976 1216
rect 364616 1164 364668 1216
rect 366548 1164 366600 1216
rect 371332 1164 371384 1216
rect 378692 1164 378744 1216
rect 384396 1164 384448 1216
rect 387524 1164 387576 1216
rect 394240 1164 394292 1216
rect 395252 1164 395304 1216
rect 402520 1164 402572 1216
rect 412916 1164 412968 1216
rect 421380 1164 421432 1216
rect 421748 1164 421800 1216
rect 430856 1164 430908 1216
rect 439412 1164 439464 1216
rect 443552 1164 443604 1216
rect 445852 1232 445904 1284
rect 449348 1232 449400 1284
rect 456984 1300 457036 1352
rect 457076 1300 457128 1352
rect 468300 1300 468352 1352
rect 481364 1300 481416 1352
rect 494704 1300 494756 1352
rect 495716 1300 495768 1352
rect 509700 1300 509752 1352
rect 510068 1300 510120 1352
rect 525432 1300 525484 1352
rect 539876 1300 539928 1352
rect 556988 1300 557040 1352
rect 454868 1232 454920 1284
rect 448612 1164 448664 1216
rect 450452 1164 450504 1216
rect 462596 1232 462648 1284
rect 474188 1232 474240 1284
rect 480168 1232 480220 1284
rect 493140 1232 493192 1284
rect 493508 1232 493560 1284
rect 507308 1232 507360 1284
rect 507768 1232 507820 1284
rect 517520 1232 517572 1284
rect 534356 1232 534408 1284
rect 551100 1232 551152 1284
rect 352196 1096 352248 1148
rect 356336 1096 356388 1148
rect 361028 1096 361080 1148
rect 365444 1096 365496 1148
rect 367652 1096 367704 1148
rect 372896 1096 372948 1148
rect 375288 1096 375340 1148
rect 4068 1028 4120 1080
rect 23112 1028 23164 1080
rect 355508 1028 355560 1080
rect 359924 1028 359976 1080
rect 373172 1028 373224 1080
rect 378508 1028 378560 1080
rect 379796 1096 379848 1148
rect 385960 1096 386012 1148
rect 386328 1096 386380 1148
rect 392676 1096 392728 1148
rect 397368 1096 397420 1148
rect 404820 1096 404872 1148
rect 420644 1096 420696 1148
rect 429292 1096 429344 1148
rect 434996 1096 435048 1148
rect 445024 1096 445076 1148
rect 445208 1096 445260 1148
rect 455696 1096 455748 1148
rect 465908 1164 465960 1216
rect 475844 1164 475896 1216
rect 488816 1164 488868 1216
rect 501236 1164 501288 1216
rect 515496 1164 515548 1216
rect 516692 1164 516744 1216
rect 532056 1164 532108 1216
rect 461584 1096 461636 1148
rect 469128 1096 469180 1148
rect 481364 1096 481416 1148
rect 487988 1096 488040 1148
rect 501420 1096 501472 1148
rect 506756 1096 506808 1148
rect 517612 1096 517664 1148
rect 522212 1096 522264 1148
rect 538128 1096 538180 1148
rect 381176 1028 381228 1080
rect 385316 1028 385368 1080
rect 391848 1028 391900 1080
rect 394148 1028 394200 1080
rect 401324 1028 401376 1080
rect 415124 1028 415176 1080
rect 423404 1028 423456 1080
rect 424968 1028 425020 1080
rect 434076 1028 434128 1080
rect 441528 1028 441580 1080
rect 451740 1028 451792 1080
rect 455972 1028 456024 1080
rect 467472 1028 467524 1080
rect 474648 1028 474700 1080
rect 487252 1028 487304 1080
rect 518808 1028 518860 1080
rect 534540 1028 534592 1080
rect 20628 960 20680 1012
rect 38568 960 38620 1012
rect 345572 960 345624 1012
rect 349252 960 349304 1012
rect 351092 960 351144 1012
rect 355232 960 355284 1012
rect 362132 960 362184 1012
rect 367008 960 367060 1012
rect 369768 960 369820 1012
rect 375288 960 375340 1012
rect 376484 960 376536 1012
rect 382372 960 382424 1012
rect 422852 960 422904 1012
rect 431868 960 431920 1012
rect 432788 960 432840 1012
rect 442632 960 442684 1012
rect 443552 960 443604 1012
rect 449808 960 449860 1012
rect 489092 960 489144 1012
rect 502984 960 503036 1012
rect 520004 960 520056 1012
rect 536104 960 536156 1012
rect 1676 892 1728 944
rect 20904 892 20956 944
rect 358728 892 358780 944
rect 363512 892 363564 944
rect 416228 892 416280 944
rect 424968 892 425020 944
rect 433892 892 433944 944
rect 443460 892 443512 944
rect 446036 892 446088 944
rect 456892 892 456944 944
rect 494612 892 494664 944
rect 508872 892 508924 944
rect 515588 892 515640 944
rect 525800 892 525852 944
rect 532148 892 532200 944
rect 548708 892 548760 944
rect 19432 824 19484 876
rect 37464 824 37516 876
rect 337844 824 337896 876
rect 340972 824 341024 876
rect 347688 824 347740 876
rect 351644 824 351696 876
rect 368756 824 368808 876
rect 373908 824 373960 876
rect 448244 824 448296 876
rect 459192 824 459244 876
rect 485688 824 485740 876
rect 498936 824 498988 876
rect 527732 824 527784 876
rect 544384 824 544436 876
rect 547604 824 547656 876
rect 565636 824 565688 876
rect 18236 756 18288 808
rect 36360 756 36412 808
rect 251180 756 251232 808
rect 253848 756 253900 808
rect 427268 756 427320 808
rect 436744 756 436796 808
rect 442724 756 442776 808
rect 453304 756 453356 808
rect 9956 688 10008 740
rect 28632 688 28684 740
rect 401876 688 401928 740
rect 409236 688 409288 740
rect 429476 688 429528 740
rect 439136 688 439188 740
rect 440516 688 440568 740
rect 450912 688 450964 740
rect 451556 688 451608 740
rect 462412 756 462464 808
rect 483572 756 483624 808
rect 497096 756 497148 808
rect 499028 756 499080 808
rect 513564 756 513616 808
rect 528836 756 528888 808
rect 545488 756 545540 808
rect 550916 756 550968 808
rect 569132 756 569184 808
rect 468116 688 468168 740
rect 480536 688 480588 740
rect 482468 688 482520 740
rect 495532 688 495584 740
rect 502248 688 502300 740
rect 517152 688 517204 740
rect 521108 688 521160 740
rect 537208 688 537260 740
rect 537668 688 537720 740
rect 554964 688 555016 740
rect 8760 620 8812 672
rect 27528 620 27580 672
rect 34796 620 34848 672
rect 51816 620 51868 672
rect 393044 620 393096 672
rect 400128 620 400180 672
rect 400772 620 400824 672
rect 408592 620 408644 672
rect 409604 620 409656 672
rect 417884 620 417936 672
rect 14740 552 14792 604
rect 17040 552 17092 604
rect 35256 552 35308 604
rect 35992 552 36044 604
rect 52920 552 52972 604
rect 389732 552 389784 604
rect 396540 552 396592 604
rect 408408 552 408460 604
rect 416688 552 416740 604
rect 431684 552 431736 604
rect 441528 620 441580 672
rect 456984 620 457036 672
rect 460020 620 460072 672
rect 464804 620 464856 672
rect 476948 620 477000 672
rect 486884 620 486936 672
rect 500592 620 500644 672
rect 503444 620 503496 672
rect 518348 620 518400 672
rect 523316 620 523368 672
rect 33048 484 33100 536
rect 39764 484 39816 536
rect 56232 484 56284 536
rect 430488 484 430540 536
rect 440332 552 440384 604
rect 447048 552 447100 604
rect 458088 552 458140 604
rect 461492 552 461544 604
rect 473452 552 473504 604
rect 486424 552 486476 604
rect 459468 484 459520 536
rect 470784 484 470836 536
rect 473636 484 473688 536
rect 16212 416 16264 468
rect 34152 416 34204 468
rect 38568 416 38620 468
rect 55128 416 55180 468
rect 382004 416 382056 468
rect 387892 416 387944 468
rect 412088 416 412140 468
rect 420368 416 420420 468
rect 437204 416 437256 468
rect 447232 416 447284 468
rect 470324 416 470376 468
rect 482468 416 482520 468
rect 484676 416 484728 468
rect 498200 552 498252 604
rect 490196 416 490248 468
rect 503812 552 503864 604
rect 508964 552 509016 604
rect 523868 552 523920 604
rect 524328 620 524380 672
rect 533252 620 533304 672
rect 539600 620 539652 672
rect 542084 620 542136 672
rect 533712 552 533764 604
rect 533804 552 533856 604
rect 11520 348 11572 400
rect 29736 348 29788 400
rect 32220 348 32272 400
rect 49608 348 49660 400
rect 407396 348 407448 400
rect 415308 348 415360 400
rect 460572 348 460624 400
rect 472440 348 472492 400
rect 478328 348 478380 400
rect 490748 348 490800 400
rect 497924 348 497976 400
rect 512092 484 512144 536
rect 517796 484 517848 536
rect 500132 416 500184 468
rect 514944 416 514996 468
rect 525708 416 525760 468
rect 542176 416 542228 468
rect 504548 348 504600 400
rect 519728 348 519780 400
rect 533252 348 533304 400
rect 540428 348 540480 400
rect 548984 620 549036 672
rect 566832 620 566884 672
rect 545396 552 545448 604
rect 563244 552 563296 604
rect 559380 484 559432 536
rect 544568 416 544620 468
rect 562232 416 562284 468
rect 550456 348 550508 400
rect 555332 348 555384 400
rect 573548 348 573600 400
rect 3240 280 3292 332
rect 22008 280 22060 332
rect 30288 280 30340 332
rect 47400 280 47452 332
rect 398564 280 398616 332
rect 406200 280 406252 332
rect 410984 280 411036 332
rect 418620 280 418672 332
rect 453764 280 453816 332
rect 464988 280 465040 332
rect 471428 280 471480 332
rect 484216 280 484268 332
rect 505652 280 505704 332
rect 520372 280 520424 332
rect 531044 280 531096 332
rect 548064 280 548116 332
rect 551928 280 551980 332
rect 570512 280 570564 332
rect 22836 212 22888 264
rect 40500 212 40552 264
rect 42248 212 42300 264
rect 58164 212 58216 264
rect 354404 212 354456 264
rect 358912 212 358964 264
rect 380808 212 380860 264
rect 386788 212 386840 264
rect 391664 212 391716 264
rect 398748 212 398800 264
rect 405188 212 405240 264
rect 412824 212 412876 264
rect 457904 212 457956 264
rect 470048 212 470100 264
rect 472532 212 472584 264
rect 484860 212 484912 264
rect 511448 212 511500 264
rect 526260 212 526312 264
rect 538772 212 538824 264
rect 556344 212 556396 264
rect 557172 212 557224 264
rect 575940 212 575992 264
rect 8024 144 8076 196
rect 26332 144 26384 196
rect 31116 144 31168 196
rect 48504 144 48556 196
rect 53564 144 53616 196
rect 69480 144 69532 196
rect 418436 144 418488 196
rect 426900 144 426952 196
rect 465816 144 465868 196
rect 478328 144 478380 196
rect 479156 144 479208 196
rect 492496 144 492548 196
rect 492588 144 492640 196
rect 506664 144 506716 196
rect 512644 144 512696 196
rect 528008 144 528060 196
rect 535368 144 535420 196
rect 552848 144 552900 196
rect 554228 144 554280 196
rect 572904 144 572956 196
rect 22008 76 22060 128
rect 39396 76 39448 128
rect 45284 76 45336 128
rect 61752 76 61804 128
rect 399668 76 399720 128
rect 407028 76 407080 128
rect 423956 76 424008 128
rect 433432 76 433484 128
rect 452568 76 452620 128
rect 464160 76 464212 128
rect 467012 76 467064 128
rect 478972 76 479024 128
rect 491300 76 491352 128
rect 505560 76 505612 128
rect 514484 76 514536 128
rect 529940 76 529992 128
rect 540980 76 541032 128
rect 558736 76 558788 128
rect 558828 76 558880 128
rect 577136 76 577188 128
rect 388 8 440 60
rect 19800 8 19852 60
rect 24584 8 24636 60
rect 41604 8 41656 60
rect 42892 8 42944 60
rect 59360 8 59412 60
rect 344744 8 344796 60
rect 348240 8 348292 60
rect 363236 8 363288 60
rect 367836 8 367888 60
rect 383108 8 383160 60
rect 389640 8 389692 60
rect 390836 8 390888 60
rect 397920 8 397972 60
rect 402888 8 402940 60
rect 410984 8 411036 60
rect 417332 8 417384 60
rect 425796 8 425848 60
rect 463608 8 463660 60
rect 475936 8 475988 60
rect 477224 8 477276 60
rect 490104 8 490156 60
rect 496728 8 496780 60
rect 511448 8 511500 60
rect 526904 8 526956 60
rect 542820 8 542872 60
rect 546408 8 546460 60
rect 564624 8 564676 60
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 251652 703582 251864 703610
rect 8128 701010 8156 703520
rect 24320 702506 24348 703520
rect 24308 702500 24360 702506
rect 24308 702442 24360 702448
rect 29276 702500 29328 702506
rect 29276 702442 29328 702448
rect 8116 701004 8168 701010
rect 8116 700946 8168 700952
rect 13084 701004 13136 701010
rect 13084 700946 13136 700952
rect 13096 700890 13124 700946
rect 13096 700862 13386 700890
rect 29288 700876 29316 702442
rect 40512 701010 40540 703520
rect 56796 701010 56824 703520
rect 72988 701010 73016 703520
rect 89180 701010 89208 703520
rect 105464 701010 105492 703520
rect 121656 701010 121684 703520
rect 137848 701010 137876 703520
rect 154132 701010 154160 703520
rect 170324 701010 170352 703520
rect 186516 703050 186544 703520
rect 186504 703044 186556 703050
rect 186504 702986 186556 702992
rect 188436 703044 188488 703050
rect 188436 702986 188488 702992
rect 40500 701004 40552 701010
rect 40500 700946 40552 700952
rect 44916 701004 44968 701010
rect 44916 700946 44968 700952
rect 56784 701004 56836 701010
rect 56784 700946 56836 700952
rect 60740 701004 60792 701010
rect 60740 700946 60792 700952
rect 72976 701004 73028 701010
rect 72976 700946 73028 700952
rect 76748 701004 76800 701010
rect 76748 700946 76800 700952
rect 89168 701004 89220 701010
rect 89168 700946 89220 700952
rect 92572 701004 92624 701010
rect 92572 700946 92624 700952
rect 105452 701004 105504 701010
rect 105452 700946 105504 700952
rect 108580 701004 108632 701010
rect 108580 700946 108632 700952
rect 121644 701004 121696 701010
rect 121644 700946 121696 700952
rect 124404 701004 124456 701010
rect 124404 700946 124456 700952
rect 137836 701004 137888 701010
rect 137836 700946 137888 700952
rect 140412 701004 140464 701010
rect 140412 700946 140464 700952
rect 154120 701004 154172 701010
rect 154120 700946 154172 700952
rect 156236 701004 156288 701010
rect 156236 700946 156288 700952
rect 170312 701004 170364 701010
rect 170312 700946 170364 700952
rect 172428 701004 172480 701010
rect 172428 700946 172480 700952
rect 44928 700890 44956 700946
rect 60752 700890 60780 700946
rect 76760 700890 76788 700946
rect 92584 700890 92612 700946
rect 108592 700890 108620 700946
rect 124416 700890 124444 700946
rect 140424 700890 140452 700946
rect 156248 700890 156276 700946
rect 172440 700890 172468 700946
rect 44928 700862 45218 700890
rect 60752 700862 61134 700890
rect 76760 700862 77050 700890
rect 92584 700862 92966 700890
rect 108592 700862 108882 700890
rect 124416 700862 124798 700890
rect 140424 700862 140714 700890
rect 156248 700862 156630 700890
rect 172440 700862 172546 700890
rect 188448 700876 188476 702986
rect 202800 701010 202828 703520
rect 218992 702506 219020 703520
rect 235184 703050 235212 703520
rect 251468 703474 251496 703520
rect 251652 703474 251680 703582
rect 251468 703446 251680 703474
rect 235172 703044 235224 703050
rect 235172 702986 235224 702992
rect 236184 703044 236236 703050
rect 236184 702986 236236 702992
rect 218980 702500 219032 702506
rect 218980 702442 219032 702448
rect 220268 702500 220320 702506
rect 220268 702442 220320 702448
rect 202788 701004 202840 701010
rect 202788 700946 202840 700952
rect 204260 701004 204312 701010
rect 204260 700946 204312 700952
rect 204272 700890 204300 700946
rect 204272 700862 204378 700890
rect 220280 700876 220308 702442
rect 236196 700876 236224 702986
rect 251836 700890 251864 703582
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332152 703582 332364 703610
rect 267660 700890 267688 703520
rect 283852 700890 283880 703520
rect 300136 700890 300164 703520
rect 316328 702434 316356 703520
rect 316052 702406 316356 702434
rect 316052 700890 316080 702406
rect 332152 700890 332180 703582
rect 332336 703474 332364 703582
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 332520 703474 332548 703520
rect 332336 703446 332548 703474
rect 348804 701010 348832 703520
rect 364996 701010 365024 703520
rect 381188 701010 381216 703520
rect 397472 701010 397500 703520
rect 413664 701010 413692 703520
rect 429856 701010 429884 703520
rect 446140 701010 446168 703520
rect 462332 702506 462360 703520
rect 459100 702500 459152 702506
rect 459100 702442 459152 702448
rect 462320 702500 462372 702506
rect 462320 702442 462372 702448
rect 348056 701004 348108 701010
rect 348056 700946 348108 700952
rect 348792 701004 348844 701010
rect 348792 700946 348844 700952
rect 363880 701004 363932 701010
rect 363880 700946 363932 700952
rect 364984 701004 365036 701010
rect 364984 700946 365036 700952
rect 379336 701004 379388 701010
rect 379336 700946 379388 700952
rect 381176 701004 381228 701010
rect 381176 700946 381228 700952
rect 395712 701004 395764 701010
rect 395712 700946 395764 700952
rect 397460 701004 397512 701010
rect 397460 700946 397512 700952
rect 411720 701004 411772 701010
rect 411720 700946 411772 700952
rect 413652 701004 413704 701010
rect 413652 700946 413704 700952
rect 427544 701004 427596 701010
rect 427544 700946 427596 700952
rect 429844 701004 429896 701010
rect 429844 700946 429896 700952
rect 443552 701004 443604 701010
rect 443552 700946 443604 700952
rect 446128 701004 446180 701010
rect 446128 700946 446180 700952
rect 348068 700890 348096 700946
rect 363892 700890 363920 700946
rect 251836 700862 252126 700890
rect 267660 700862 268042 700890
rect 283852 700862 283958 700890
rect 299966 700862 300164 700890
rect 315882 700862 316080 700890
rect 331798 700862 332180 700890
rect 347714 700862 348096 700890
rect 363630 700862 363920 700890
rect 379348 700890 379376 700946
rect 395724 700890 395752 700946
rect 411732 700890 411760 700946
rect 427556 700890 427584 700946
rect 443564 700890 443592 700946
rect 379348 700862 379454 700890
rect 395462 700862 395752 700890
rect 411378 700862 411760 700890
rect 427294 700862 427584 700890
rect 443210 700862 443592 700890
rect 459112 700876 459140 702442
rect 478524 701010 478552 703520
rect 494808 702778 494836 703520
rect 490932 702772 490984 702778
rect 490932 702714 490984 702720
rect 494796 702772 494848 702778
rect 494796 702714 494848 702720
rect 475384 701004 475436 701010
rect 475384 700946 475436 700952
rect 478512 701004 478564 701010
rect 478512 700946 478564 700952
rect 475396 700890 475424 700946
rect 475042 700862 475424 700890
rect 490944 700876 490972 702714
rect 511000 702506 511028 703520
rect 527192 703066 527220 703520
rect 527100 703050 527220 703066
rect 522764 703044 522816 703050
rect 522764 702986 522816 702992
rect 527088 703044 527220 703050
rect 527140 703038 527220 703044
rect 527088 702986 527140 702992
rect 506848 702500 506900 702506
rect 506848 702442 506900 702448
rect 510988 702500 511040 702506
rect 510988 702442 511040 702448
rect 506860 700876 506888 702442
rect 522776 700876 522804 702986
rect 543476 702778 543504 703520
rect 538680 702772 538732 702778
rect 538680 702714 538732 702720
rect 543464 702772 543516 702778
rect 543464 702714 543516 702720
rect 538692 700876 538720 702714
rect 559668 702506 559696 703520
rect 575860 703050 575888 703520
rect 570512 703044 570564 703050
rect 570512 702986 570564 702992
rect 575848 703044 575900 703050
rect 575848 702986 575900 702992
rect 554596 702500 554648 702506
rect 554596 702442 554648 702448
rect 559656 702500 559708 702506
rect 559656 702442 559708 702448
rect 554608 700876 554636 702442
rect 570524 700876 570552 702986
rect 2778 697368 2834 697377
rect 2778 697303 2834 697312
rect 2792 690849 2820 697303
rect 581642 697232 581698 697241
rect 581642 697167 581698 697176
rect 581656 691529 581684 697167
rect 581642 691520 581698 691529
rect 581642 691455 581698 691464
rect 2778 690840 2834 690849
rect 2778 690775 2834 690784
rect 2778 684312 2834 684321
rect 2778 684247 2834 684256
rect 2792 678065 2820 684247
rect 582378 683904 582434 683913
rect 582378 683839 582434 683848
rect 582392 678473 582420 683839
rect 582378 678464 582434 678473
rect 582378 678399 582434 678408
rect 2778 678056 2834 678065
rect 2778 677991 2834 678000
rect 2778 671256 2834 671265
rect 2778 671191 2834 671200
rect 2792 665281 2820 671191
rect 582378 670712 582434 670721
rect 582378 670647 582434 670656
rect 582392 665417 582420 670647
rect 582378 665408 582434 665417
rect 582378 665343 582434 665352
rect 2778 665272 2834 665281
rect 2778 665207 2834 665216
rect 2778 658200 2834 658209
rect 2778 658135 2834 658144
rect 2792 652497 2820 658135
rect 582378 657384 582434 657393
rect 582378 657319 582434 657328
rect 2778 652488 2834 652497
rect 2778 652423 2834 652432
rect 582392 652361 582420 657319
rect 582378 652352 582434 652361
rect 582378 652287 582434 652296
rect 2778 645144 2834 645153
rect 2778 645079 2834 645088
rect 2792 639713 2820 645079
rect 581642 644056 581698 644065
rect 581642 643991 581698 644000
rect 2778 639704 2834 639713
rect 2778 639639 2834 639648
rect 581656 639305 581684 643991
rect 581642 639296 581698 639305
rect 581642 639231 581698 639240
rect 2778 632088 2834 632097
rect 2778 632023 2834 632032
rect 2792 626929 2820 632023
rect 582378 630864 582434 630873
rect 582378 630799 582434 630808
rect 2778 626920 2834 626929
rect 2778 626855 2834 626864
rect 582392 626249 582420 630799
rect 582378 626240 582434 626249
rect 582378 626175 582434 626184
rect 2778 619168 2834 619177
rect 2778 619103 2834 619112
rect 2792 614009 2820 619103
rect 581642 617536 581698 617545
rect 581642 617471 581698 617480
rect 2778 614000 2834 614009
rect 2778 613935 2834 613944
rect 581656 613193 581684 617471
rect 581642 613184 581698 613193
rect 581642 613119 581698 613128
rect 2778 606112 2834 606121
rect 2778 606047 2834 606056
rect 2792 601361 2820 606047
rect 581642 604208 581698 604217
rect 581642 604143 581698 604152
rect 2778 601352 2834 601361
rect 2778 601287 2834 601296
rect 581656 600137 581684 604143
rect 581642 600128 581698 600137
rect 581642 600063 581698 600072
rect 1582 593056 1638 593065
rect 1582 592991 1638 593000
rect 1596 588577 1624 592991
rect 581642 591016 581698 591025
rect 581642 590951 581698 590960
rect 1582 588568 1638 588577
rect 1582 588503 1638 588512
rect 581656 587081 581684 590951
rect 581642 587072 581698 587081
rect 581642 587007 581698 587016
rect 2042 580000 2098 580009
rect 2042 579935 2098 579944
rect 2056 575793 2084 579935
rect 581642 577688 581698 577697
rect 581642 577623 581698 577632
rect 2042 575784 2098 575793
rect 2042 575719 2098 575728
rect 581656 574025 581684 577623
rect 581642 574016 581698 574025
rect 581642 573951 581698 573960
rect 1490 566944 1546 566953
rect 1490 566879 1546 566888
rect 1504 563009 1532 566879
rect 582378 564360 582434 564369
rect 582378 564295 582434 564304
rect 1490 563000 1546 563009
rect 1490 562935 1546 562944
rect 582392 560969 582420 564295
rect 582378 560960 582434 560969
rect 582378 560895 582434 560904
rect 1490 553888 1546 553897
rect 1490 553823 1546 553832
rect 1504 550225 1532 553823
rect 581642 551168 581698 551177
rect 581642 551103 581698 551112
rect 1490 550216 1546 550225
rect 1490 550151 1546 550160
rect 581656 547777 581684 551103
rect 581642 547768 581698 547777
rect 581642 547703 581698 547712
rect 1398 540832 1454 540841
rect 1398 540767 1454 540776
rect 1412 537441 1440 540767
rect 582378 537840 582434 537849
rect 582378 537775 582434 537784
rect 1398 537432 1454 537441
rect 1398 537367 1454 537376
rect 582392 534857 582420 537775
rect 582378 534848 582434 534857
rect 582378 534783 582434 534792
rect 1490 527912 1546 527921
rect 1490 527847 1546 527856
rect 1504 524657 1532 527847
rect 1490 524648 1546 524657
rect 1490 524583 1546 524592
rect 582378 524512 582434 524521
rect 582378 524447 582434 524456
rect 582392 521801 582420 524447
rect 582378 521792 582434 521801
rect 582378 521727 582434 521736
rect 1582 514856 1638 514865
rect 1582 514791 1638 514800
rect 1596 511873 1624 514791
rect 1582 511864 1638 511873
rect 1582 511799 1638 511808
rect 582378 511320 582434 511329
rect 582378 511255 582434 511264
rect 582392 508745 582420 511255
rect 582378 508736 582434 508745
rect 582378 508671 582434 508680
rect 1582 501800 1638 501809
rect 1582 501735 1638 501744
rect 1596 499089 1624 501735
rect 1582 499080 1638 499089
rect 1582 499015 1638 499024
rect 581642 497992 581698 498001
rect 581642 497927 581698 497936
rect 581656 495689 581684 497927
rect 581642 495680 581698 495689
rect 581642 495615 581698 495624
rect 1582 488744 1638 488753
rect 1582 488679 1638 488688
rect 1596 486305 1624 488679
rect 1582 486296 1638 486305
rect 1582 486231 1638 486240
rect 582378 484664 582434 484673
rect 582378 484599 582434 484608
rect 582392 482633 582420 484599
rect 582378 482624 582434 482633
rect 582378 482559 582434 482568
rect 2778 475688 2834 475697
rect 2778 475623 2834 475632
rect 2792 473521 2820 475623
rect 2778 473512 2834 473521
rect 2778 473447 2834 473456
rect 581642 471472 581698 471481
rect 581642 471407 581698 471416
rect 581656 469577 581684 471407
rect 581642 469568 581698 469577
rect 581642 469503 581698 469512
rect 1582 462632 1638 462641
rect 1582 462567 1638 462576
rect 1596 460737 1624 462567
rect 1582 460728 1638 460737
rect 1582 460663 1638 460672
rect 581642 458144 581698 458153
rect 581642 458079 581698 458088
rect 581656 456521 581684 458079
rect 581642 456512 581698 456521
rect 581642 456447 581698 456456
rect 2778 449576 2834 449585
rect 2778 449511 2834 449520
rect 2792 447953 2820 449511
rect 2778 447944 2834 447953
rect 2778 447879 2834 447888
rect 2778 436656 2834 436665
rect 2778 436591 2834 436600
rect 2792 435169 2820 436591
rect 2778 435160 2834 435169
rect 2778 435095 2834 435104
rect 2778 423600 2834 423609
rect 2778 423535 2834 423544
rect 2792 422385 2820 423535
rect 2778 422376 2834 422385
rect 2778 422311 2834 422320
rect 1306 294400 1362 294409
rect 1306 294335 1362 294344
rect 1320 293185 1348 294335
rect 1306 293176 1362 293185
rect 1306 293111 1362 293120
rect 2778 281616 2834 281625
rect 2778 281551 2834 281560
rect 2792 280129 2820 281551
rect 2778 280120 2834 280129
rect 2778 280055 2834 280064
rect 1306 268832 1362 268841
rect 1306 268767 1362 268776
rect 1320 267209 1348 268767
rect 1306 267200 1362 267209
rect 1306 267135 1362 267144
rect 582378 260536 582434 260545
rect 582378 260471 582434 260480
rect 582392 258913 582420 260471
rect 582378 258904 582434 258913
rect 582378 258839 582434 258848
rect 1306 256048 1362 256057
rect 1306 255983 1362 255992
rect 1320 254153 1348 255983
rect 1306 254144 1362 254153
rect 1306 254079 1362 254088
rect 580906 247072 580962 247081
rect 580906 247007 580962 247016
rect 580920 245585 580948 247007
rect 580906 245576 580962 245585
rect 580906 245511 580962 245520
rect 2778 243264 2834 243273
rect 2778 243199 2834 243208
rect 2792 241097 2820 243199
rect 2778 241088 2834 241097
rect 2778 241023 2834 241032
rect 582378 234424 582434 234433
rect 582378 234359 582434 234368
rect 582392 232393 582420 234359
rect 582378 232384 582434 232393
rect 582378 232319 582434 232328
rect 2778 230616 2834 230625
rect 2778 230551 2834 230560
rect 2792 228041 2820 230551
rect 2778 228032 2834 228041
rect 2778 227967 2834 227976
rect 580906 220960 580962 220969
rect 580906 220895 580962 220904
rect 580920 219065 580948 220895
rect 580906 219056 580962 219065
rect 580906 218991 580962 219000
rect 2778 217696 2834 217705
rect 2778 217631 2834 217640
rect 2792 214985 2820 217631
rect 2778 214976 2834 214985
rect 2778 214911 2834 214920
rect 582378 208312 582434 208321
rect 582378 208247 582434 208256
rect 582392 205737 582420 208247
rect 582378 205728 582434 205737
rect 582378 205663 582434 205672
rect 2778 204912 2834 204921
rect 2778 204847 2834 204856
rect 2792 201929 2820 204847
rect 2778 201920 2834 201929
rect 2778 201855 2834 201864
rect 580906 194712 580962 194721
rect 580906 194647 580962 194656
rect 580920 192545 580948 194647
rect 580906 192536 580962 192545
rect 580906 192471 580962 192480
rect 1306 192128 1362 192137
rect 1306 192063 1362 192072
rect 1320 188873 1348 192063
rect 1306 188864 1362 188873
rect 1306 188799 1362 188808
rect 580906 182472 580962 182481
rect 580906 182407 580962 182416
rect 2778 179344 2834 179353
rect 2778 179279 2834 179288
rect 2792 175953 2820 179279
rect 580920 179217 580948 182407
rect 580906 179208 580962 179217
rect 580906 179143 580962 179152
rect 2778 175944 2834 175953
rect 2778 175879 2834 175888
rect 580906 168600 580962 168609
rect 580906 168535 580962 168544
rect 2778 166560 2834 166569
rect 2778 166495 2834 166504
rect 2792 162897 2820 166495
rect 580920 165889 580948 168535
rect 580906 165880 580962 165889
rect 580906 165815 580962 165824
rect 2778 162888 2834 162897
rect 2778 162823 2834 162832
rect 580906 156360 580962 156369
rect 580906 156295 580962 156304
rect 1306 153776 1362 153785
rect 1306 153711 1362 153720
rect 1320 149841 1348 153711
rect 580920 152697 580948 156295
rect 580906 152688 580962 152697
rect 580906 152623 580962 152632
rect 1306 149832 1362 149841
rect 1306 149767 1362 149776
rect 580906 142624 580962 142633
rect 580906 142559 580962 142568
rect 570 140992 626 141001
rect 570 140927 626 140936
rect 584 136785 612 140927
rect 580920 139369 580948 142559
rect 580906 139360 580962 139369
rect 580906 139295 580962 139304
rect 570 136776 626 136785
rect 570 136711 626 136720
rect 580906 130248 580962 130257
rect 580906 130183 580962 130192
rect 754 128208 810 128217
rect 754 128143 810 128152
rect 768 123729 796 128143
rect 580920 126041 580948 130183
rect 580906 126032 580962 126041
rect 580906 125967 580962 125976
rect 754 123720 810 123729
rect 754 123655 810 123664
rect 579894 116376 579950 116385
rect 579894 116311 579950 116320
rect 1306 115424 1362 115433
rect 1306 115359 1362 115368
rect 1320 110673 1348 115359
rect 579908 112849 579936 116311
rect 579894 112840 579950 112849
rect 579894 112775 579950 112784
rect 1306 110664 1362 110673
rect 1306 110599 1362 110608
rect 580906 103592 580962 103601
rect 580906 103527 580962 103536
rect 1582 102640 1638 102649
rect 1582 102575 1638 102584
rect 1596 97617 1624 102575
rect 580920 99521 580948 103527
rect 580906 99512 580962 99521
rect 580906 99447 580962 99456
rect 1582 97608 1638 97617
rect 1582 97543 1638 97552
rect 580906 90264 580962 90273
rect 580906 90199 580962 90208
rect 1582 89856 1638 89865
rect 1582 89791 1638 89800
rect 1596 84697 1624 89791
rect 580920 86193 580948 90199
rect 580906 86184 580962 86193
rect 580906 86119 580962 86128
rect 1582 84688 1638 84697
rect 1582 84623 1638 84632
rect 579894 77344 579950 77353
rect 579894 77279 579950 77288
rect 1582 77072 1638 77081
rect 1582 77007 1638 77016
rect 1596 71641 1624 77007
rect 579908 73001 579936 77279
rect 579894 72992 579950 73001
rect 579894 72927 579950 72936
rect 1582 71632 1638 71641
rect 1582 71567 1638 71576
rect 1490 64288 1546 64297
rect 1490 64223 1546 64232
rect 1504 58585 1532 64223
rect 580906 64152 580962 64161
rect 580906 64087 580962 64096
rect 580920 59673 580948 64087
rect 580906 59664 580962 59673
rect 580906 59599 580962 59608
rect 1490 58576 1546 58585
rect 1490 58511 1546 58520
rect 2042 51504 2098 51513
rect 2042 51439 2098 51448
rect 2056 45529 2084 51439
rect 580906 51096 580962 51105
rect 580906 51031 580962 51040
rect 580920 46345 580948 51031
rect 580906 46336 580962 46345
rect 580906 46271 580962 46280
rect 2042 45520 2098 45529
rect 2042 45455 2098 45464
rect 2042 38720 2098 38729
rect 2042 38655 2098 38664
rect 2056 32473 2084 38655
rect 580906 38040 580962 38049
rect 580906 37975 580962 37984
rect 580920 33153 580948 37975
rect 580906 33144 580962 33153
rect 580906 33079 580962 33088
rect 2042 32464 2098 32473
rect 2042 32399 2098 32408
rect 1490 25936 1546 25945
rect 1490 25871 1546 25880
rect 1504 19417 1532 25871
rect 580906 24984 580962 24993
rect 580906 24919 580962 24928
rect 580920 19825 580948 24919
rect 580906 19816 580962 19825
rect 580906 19751 580962 19760
rect 1490 19408 1546 19417
rect 1490 19343 1546 19352
rect 2042 13152 2098 13161
rect 2042 13087 2098 13096
rect 2056 6497 2084 13087
rect 579894 12744 579950 12753
rect 579894 12679 579950 12688
rect 579908 6633 579936 12679
rect 579894 6624 579950 6633
rect 579894 6559 579950 6568
rect 2042 6488 2098 6497
rect 2042 6423 2098 6432
rect 74736 4010 75026 4026
rect 74724 4004 75026 4010
rect 74776 3998 75026 4004
rect 74724 3946 74776 3952
rect 70216 3936 70268 3942
rect 70214 3904 70216 3913
rect 78036 3936 78088 3942
rect 70268 3904 70270 3913
rect 59728 3868 59780 3874
rect 70214 3839 70270 3848
rect 73618 3904 73674 3913
rect 73674 3862 73922 3890
rect 78088 3884 78338 3890
rect 78036 3878 78338 3884
rect 78048 3862 78338 3878
rect 83568 3874 83858 3890
rect 94608 3874 94898 3890
rect 133248 3874 133538 3890
rect 83556 3868 83858 3874
rect 73618 3839 73674 3848
rect 59728 3810 59780 3816
rect 83608 3862 83858 3868
rect 94596 3868 94898 3874
rect 83556 3810 83608 3816
rect 94648 3862 94898 3868
rect 122288 3868 122340 3874
rect 94596 3810 94648 3816
rect 122288 3810 122340 3816
rect 133236 3868 133538 3874
rect 133288 3862 133538 3868
rect 133236 3810 133288 3816
rect 58808 3732 58860 3738
rect 58808 3674 58860 3680
rect 56048 3528 56100 3534
rect 56048 3470 56100 3476
rect 54944 3460 54996 3466
rect 54944 3402 54996 3408
rect 51356 3392 51408 3398
rect 51356 3334 51408 3340
rect 50160 3256 50212 3262
rect 50160 3198 50212 3204
rect 40960 3188 41012 3194
rect 40960 3130 41012 3136
rect 4068 1080 4120 1086
rect 4068 1022 4120 1028
rect 1676 944 1728 950
rect 1676 886 1728 892
rect 1688 480 1716 886
rect 4080 480 4108 1022
rect 19432 876 19484 882
rect 19432 818 19484 824
rect 18236 808 18288 814
rect 18236 750 18288 756
rect 9956 740 10008 746
rect 9956 682 10008 688
rect 8760 672 8812 678
rect 8760 614 8812 620
rect 8772 480 8800 614
rect 9968 480 9996 682
rect 14740 604 14792 610
rect 14740 546 14792 552
rect 17040 604 17092 610
rect 17040 546 17092 552
rect 12162 504 12218 513
rect 542 82 654 480
rect 400 66 654 82
rect 388 60 654 66
rect 440 54 654 60
rect 388 2 440 8
rect 542 -960 654 54
rect 1646 -960 1758 480
rect 2842 354 2954 480
rect 2842 338 3280 354
rect 2842 332 3292 338
rect 2842 326 3240 332
rect 2842 -960 2954 326
rect 3240 274 3292 280
rect 4038 -960 4150 480
rect 5234 354 5346 480
rect 5446 368 5502 377
rect 5234 326 5446 354
rect 5234 -960 5346 326
rect 5446 303 5502 312
rect 6274 96 6330 105
rect 6430 82 6542 480
rect 6330 54 6542 82
rect 6274 31 6330 40
rect 6430 -960 6542 54
rect 7626 218 7738 480
rect 7626 202 8064 218
rect 7626 196 8076 202
rect 7626 190 8024 196
rect 7626 -960 7738 190
rect 8024 138 8076 144
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 354 11234 480
rect 14752 480 14780 546
rect 17052 480 17080 546
rect 18248 480 18276 750
rect 19444 480 19472 818
rect 12162 439 12218 448
rect 11520 400 11572 406
rect 11122 348 11520 354
rect 11122 342 11572 348
rect 12176 354 12204 439
rect 12318 354 12430 480
rect 11122 326 11560 342
rect 12176 326 12430 354
rect 11122 -960 11234 326
rect 12318 -960 12430 326
rect 13514 218 13626 480
rect 13726 232 13782 241
rect 13514 190 13726 218
rect 13514 -960 13626 190
rect 13726 167 13782 176
rect 14710 -960 14822 480
rect 15906 354 16018 480
rect 16212 468 16264 474
rect 16212 410 16264 416
rect 16224 354 16252 410
rect 15906 326 16252 354
rect 15906 -960 16018 326
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 19812 66 19840 3060
rect 20628 1012 20680 1018
rect 20628 954 20680 960
rect 20640 480 20668 954
rect 20916 950 20944 3060
rect 20904 944 20956 950
rect 20904 886 20956 892
rect 19800 60 19852 66
rect 19800 2 19852 8
rect 20598 -960 20710 480
rect 21794 82 21906 480
rect 22020 338 22048 3060
rect 23124 1086 23152 3060
rect 23952 3046 24242 3074
rect 25056 3046 25346 3074
rect 26344 3046 26450 3074
rect 23112 1080 23164 1086
rect 23112 1022 23164 1028
rect 22008 332 22060 338
rect 22008 274 22060 280
rect 22836 264 22888 270
rect 22990 218 23102 480
rect 23952 377 23980 3046
rect 23938 368 23994 377
rect 23938 303 23994 312
rect 22888 212 23102 218
rect 22836 206 23102 212
rect 22848 190 23102 206
rect 22008 128 22060 134
rect 21794 76 22008 82
rect 21794 70 22060 76
rect 21794 54 22048 70
rect 21794 -960 21906 54
rect 22990 -960 23102 190
rect 24186 82 24298 480
rect 25056 105 25084 3046
rect 25290 354 25402 480
rect 25686 368 25742 377
rect 25290 326 25686 354
rect 25042 96 25098 105
rect 24186 66 24624 82
rect 24186 60 24636 66
rect 24186 54 24584 60
rect 24186 -960 24298 54
rect 25042 31 25098 40
rect 24584 2 24636 8
rect 25290 -960 25402 326
rect 25686 303 25742 312
rect 26344 202 26372 3046
rect 26608 2916 26660 2922
rect 26608 2858 26660 2864
rect 26620 1442 26648 2858
rect 26528 1414 26648 1442
rect 26528 480 26556 1414
rect 27540 678 27568 3060
rect 27712 2848 27764 2854
rect 27712 2790 27764 2796
rect 27528 672 27580 678
rect 27528 614 27580 620
rect 27724 480 27752 2790
rect 28644 746 28672 3060
rect 28632 740 28684 746
rect 28632 682 28684 688
rect 28906 640 28962 649
rect 28906 575 28962 584
rect 28920 480 28948 575
rect 26332 196 26384 202
rect 26332 138 26384 144
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 29748 406 29776 3060
rect 30852 513 30880 3060
rect 30838 504 30894 513
rect 29736 400 29788 406
rect 29736 342 29788 348
rect 30074 354 30186 480
rect 30838 439 30894 448
rect 30074 338 30328 354
rect 30074 332 30340 338
rect 30074 326 30288 332
rect 30074 -960 30186 326
rect 30288 274 30340 280
rect 31270 218 31382 480
rect 31956 241 31984 3060
rect 33060 542 33088 3060
rect 33600 2984 33652 2990
rect 33600 2926 33652 2932
rect 33048 536 33100 542
rect 32220 400 32272 406
rect 32374 354 32486 480
rect 33048 478 33100 484
rect 33612 480 33640 2926
rect 32272 348 32486 354
rect 32220 342 32486 348
rect 32232 326 32486 342
rect 31128 202 31382 218
rect 31116 196 31382 202
rect 31168 190 31382 196
rect 31116 138 31168 144
rect 31270 -960 31382 190
rect 31942 232 31998 241
rect 31942 167 31998 176
rect 32374 -960 32486 326
rect 33570 -960 33682 480
rect 34164 474 34192 3060
rect 34796 672 34848 678
rect 34796 614 34848 620
rect 34808 480 34836 614
rect 35268 610 35296 3060
rect 36372 814 36400 3060
rect 37476 882 37504 3060
rect 38580 1018 38608 3060
rect 39408 3046 39698 3074
rect 40512 3046 40802 3074
rect 38568 1012 38620 1018
rect 38568 954 38620 960
rect 37464 876 37516 882
rect 37464 818 37516 824
rect 36360 808 36412 814
rect 36360 750 36412 756
rect 35256 604 35308 610
rect 35256 546 35308 552
rect 35992 604 36044 610
rect 35992 546 36044 552
rect 36004 480 36032 546
rect 34152 468 34204 474
rect 34152 410 34204 416
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37002 232 37058 241
rect 37158 218 37270 480
rect 37058 190 37270 218
rect 37002 167 37058 176
rect 37158 -960 37270 190
rect 38354 354 38466 480
rect 38568 468 38620 474
rect 38568 410 38620 416
rect 38580 354 38608 410
rect 38354 326 38608 354
rect 38354 -960 38466 326
rect 39408 134 39436 3046
rect 39592 598 39804 626
rect 39592 480 39620 598
rect 39776 542 39804 598
rect 39764 536 39816 542
rect 39396 128 39448 134
rect 39396 70 39448 76
rect 39550 -960 39662 480
rect 39764 478 39816 484
rect 40512 270 40540 3046
rect 40972 1578 41000 3130
rect 40696 1550 41000 1578
rect 41616 3046 41906 3074
rect 42812 3046 43010 3074
rect 43824 3046 44114 3074
rect 44272 3052 44324 3058
rect 40696 480 40724 1550
rect 40500 264 40552 270
rect 40500 206 40552 212
rect 40654 -960 40766 480
rect 41616 66 41644 3046
rect 41850 218 41962 480
rect 42706 368 42762 377
rect 42812 354 42840 3046
rect 43824 2922 43852 3046
rect 44272 2994 44324 3000
rect 43812 2916 43864 2922
rect 43812 2858 43864 2864
rect 44284 480 44312 2994
rect 45204 2854 45232 3060
rect 45192 2848 45244 2854
rect 45192 2790 45244 2796
rect 46308 649 46336 3060
rect 46294 640 46350 649
rect 46294 575 46350 584
rect 42762 326 42840 354
rect 42706 303 42762 312
rect 42248 264 42300 270
rect 41850 212 42248 218
rect 41850 206 42300 212
rect 41850 190 42288 206
rect 41604 60 41656 66
rect 41604 2 41656 8
rect 41850 -960 41962 190
rect 43046 82 43158 480
rect 42904 66 43158 82
rect 42892 60 43158 66
rect 42944 54 43158 60
rect 42892 2 42944 8
rect 43046 -960 43158 54
rect 44242 -960 44354 480
rect 45284 128 45336 134
rect 45438 82 45550 480
rect 45336 76 45550 82
rect 45284 70 45550 76
rect 45296 54 45550 70
rect 45438 -960 45550 54
rect 46634 82 46746 480
rect 47412 338 47440 3060
rect 47860 2848 47912 2854
rect 47860 2790 47912 2796
rect 47872 480 47900 2790
rect 47400 332 47452 338
rect 47400 274 47452 280
rect 46846 96 46902 105
rect 46634 54 46846 82
rect 46634 -960 46746 54
rect 46846 31 46902 40
rect 47830 -960 47942 480
rect 48516 202 48544 3060
rect 48964 2916 49016 2922
rect 48964 2858 49016 2864
rect 48976 480 49004 2858
rect 48504 196 48556 202
rect 48504 138 48556 144
rect 48934 -960 49046 480
rect 49620 406 49648 3060
rect 50172 480 50200 3198
rect 50448 3046 50738 3074
rect 50448 2990 50476 3046
rect 50436 2984 50488 2990
rect 50436 2926 50488 2932
rect 51368 480 51396 3334
rect 52552 3120 52604 3126
rect 52552 3062 52604 3068
rect 51828 678 51856 3060
rect 51816 672 51868 678
rect 51816 614 51868 620
rect 52564 480 52592 3062
rect 52932 610 52960 3060
rect 52920 604 52972 610
rect 52920 546 52972 552
rect 49608 400 49660 406
rect 49608 342 49660 348
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 218 53830 480
rect 54036 241 54064 3060
rect 54956 480 54984 3402
rect 53576 202 53830 218
rect 53564 196 53830 202
rect 53616 190 53830 196
rect 53564 138 53616 144
rect 53718 -960 53830 190
rect 54022 232 54078 241
rect 54022 167 54078 176
rect 54914 -960 55026 480
rect 55140 474 55168 3060
rect 56060 480 56088 3470
rect 57072 3194 57362 3210
rect 57060 3188 57362 3194
rect 57112 3182 57362 3188
rect 57520 3188 57572 3194
rect 57060 3130 57112 3136
rect 57520 3130 57572 3136
rect 56244 542 56272 3060
rect 57532 1578 57560 3130
rect 57256 1550 57560 1578
rect 58176 3046 58466 3074
rect 56232 536 56284 542
rect 55128 468 55180 474
rect 55128 410 55180 416
rect 56018 -960 56130 480
rect 56232 478 56284 484
rect 57256 480 57284 1550
rect 57214 -960 57326 480
rect 58176 270 58204 3046
rect 58410 354 58522 480
rect 58820 354 58848 3674
rect 58410 326 58848 354
rect 59372 3046 59570 3074
rect 58164 264 58216 270
rect 58164 206 58216 212
rect 58410 -960 58522 326
rect 59372 66 59400 3046
rect 59740 1986 59768 3810
rect 62028 3800 62080 3806
rect 62028 3742 62080 3748
rect 67456 3800 67508 3806
rect 80888 3800 80940 3806
rect 67456 3742 67508 3748
rect 60384 3058 60674 3074
rect 60372 3052 60674 3058
rect 60424 3046 60674 3052
rect 60372 2994 60424 3000
rect 60832 2848 60884 2854
rect 60832 2790 60884 2796
rect 59648 1958 59768 1986
rect 59648 480 59676 1958
rect 60844 480 60872 2790
rect 59360 60 59412 66
rect 59360 2 59412 8
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61764 134 61792 3060
rect 62040 480 62068 3742
rect 63224 3664 63276 3670
rect 63224 3606 63276 3612
rect 61752 128 61804 134
rect 61752 70 61804 76
rect 61998 -960 62110 480
rect 62868 105 62896 3060
rect 63236 480 63264 3606
rect 66720 3596 66772 3602
rect 66720 3538 66772 3544
rect 65524 3324 65576 3330
rect 65524 3266 65576 3272
rect 63696 3046 63986 3074
rect 64328 3052 64380 3058
rect 63696 2922 63724 3046
rect 64328 2994 64380 3000
rect 64892 3046 65090 3074
rect 63684 2916 63736 2922
rect 63684 2858 63736 2864
rect 64340 480 64368 2994
rect 64892 2990 64920 3046
rect 64880 2984 64932 2990
rect 64880 2926 64932 2932
rect 65536 480 65564 3266
rect 65892 3256 65944 3262
rect 65944 3204 66194 3210
rect 65892 3198 66194 3204
rect 65904 3182 66194 3198
rect 66732 480 66760 3538
rect 67468 3398 67496 3742
rect 71424 3738 71714 3754
rect 84476 3800 84528 3806
rect 80888 3742 80940 3748
rect 69020 3732 69072 3738
rect 69020 3674 69072 3680
rect 71412 3732 71714 3738
rect 71464 3726 71714 3732
rect 71412 3674 71464 3680
rect 69032 3534 69060 3674
rect 69112 3664 69164 3670
rect 69112 3606 69164 3612
rect 69020 3528 69072 3534
rect 69020 3470 69072 3476
rect 66996 3392 67048 3398
rect 67456 3392 67508 3398
rect 67048 3340 67298 3346
rect 66996 3334 67298 3340
rect 67456 3334 67508 3340
rect 67008 3318 67298 3334
rect 68100 3120 68152 3126
rect 68152 3068 68402 3074
rect 68100 3062 68402 3068
rect 68112 3046 68402 3062
rect 67916 2984 67968 2990
rect 67916 2926 67968 2932
rect 67928 480 67956 2926
rect 69124 480 69152 3606
rect 70124 3528 70176 3534
rect 70124 3470 70176 3476
rect 72976 3528 73028 3534
rect 72976 3470 73028 3476
rect 78588 3528 78640 3534
rect 78588 3470 78640 3476
rect 62854 96 62910 105
rect 62854 31 62910 40
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 69492 202 69520 3060
rect 70136 218 70164 3470
rect 70216 3460 70268 3466
rect 70216 3402 70268 3408
rect 70228 3346 70256 3402
rect 70228 3318 70610 3346
rect 71504 3324 71556 3330
rect 71504 3266 71556 3272
rect 71516 480 71544 3266
rect 72528 3194 72818 3210
rect 72516 3188 72818 3194
rect 72568 3182 72818 3188
rect 72516 3130 72568 3136
rect 70278 218 70390 480
rect 69480 196 69532 202
rect 70136 190 70390 218
rect 69480 138 69532 144
rect 70278 -960 70390 190
rect 71474 -960 71586 480
rect 72578 354 72690 480
rect 72988 354 73016 3470
rect 76932 3392 76984 3398
rect 76984 3340 77234 3346
rect 76932 3334 77234 3340
rect 76944 3318 77234 3334
rect 73804 3188 73856 3194
rect 73804 3130 73856 3136
rect 73816 480 73844 3130
rect 76288 3120 76340 3126
rect 75840 3046 76130 3074
rect 76288 3062 76340 3068
rect 75368 2916 75420 2922
rect 75368 2858 75420 2864
rect 72578 326 73016 354
rect 72578 -960 72690 326
rect 73774 -960 73886 480
rect 74970 354 75082 480
rect 75380 354 75408 2858
rect 75840 2854 75868 3046
rect 75828 2848 75880 2854
rect 75828 2790 75880 2796
rect 76300 1578 76328 3062
rect 77392 2848 77444 2854
rect 77392 2790 77444 2796
rect 76208 1550 76328 1578
rect 76208 480 76236 1550
rect 77404 480 77432 2790
rect 78600 480 78628 3470
rect 79692 3392 79744 3398
rect 79692 3334 79744 3340
rect 79600 3120 79652 3126
rect 79152 3058 79442 3074
rect 79600 3062 79652 3068
rect 79140 3052 79442 3058
rect 79192 3046 79442 3052
rect 79140 2994 79192 3000
rect 79612 2922 79640 3062
rect 79600 2916 79652 2922
rect 79600 2858 79652 2864
rect 79704 480 79732 3334
rect 79968 3256 80020 3262
rect 80020 3204 80546 3210
rect 79968 3198 80546 3204
rect 79980 3182 80546 3198
rect 80900 480 80928 3742
rect 81360 3738 81650 3754
rect 84476 3742 84528 3748
rect 98000 3800 98052 3806
rect 114008 3800 114060 3806
rect 98052 3748 98210 3754
rect 98000 3742 98210 3748
rect 81348 3732 81650 3738
rect 81400 3726 81650 3732
rect 81348 3674 81400 3680
rect 82912 3596 82964 3602
rect 82912 3538 82964 3544
rect 83280 3596 83332 3602
rect 83280 3538 83332 3544
rect 82924 3330 82952 3538
rect 83004 3392 83056 3398
rect 83004 3334 83056 3340
rect 82912 3324 82964 3330
rect 82912 3266 82964 3272
rect 82740 2990 82768 3060
rect 83016 3058 83044 3334
rect 83004 3052 83056 3058
rect 83004 2994 83056 3000
rect 82728 2984 82780 2990
rect 82728 2926 82780 2932
rect 82084 2916 82136 2922
rect 82084 2858 82136 2864
rect 82096 480 82124 2858
rect 83292 480 83320 3538
rect 84488 480 84516 3742
rect 85672 3732 85724 3738
rect 85672 3674 85724 3680
rect 87788 3732 87840 3738
rect 98012 3726 98210 3742
rect 101232 3738 101522 3754
rect 114008 3742 114060 3748
rect 101220 3732 101522 3738
rect 87788 3674 87840 3680
rect 101272 3726 101522 3732
rect 101220 3674 101272 3680
rect 84672 3330 84962 3346
rect 84660 3324 84962 3330
rect 84712 3318 84962 3324
rect 84660 3266 84712 3272
rect 85684 480 85712 3674
rect 86868 3664 86920 3670
rect 86920 3612 87170 3618
rect 86868 3606 87170 3612
rect 86880 3590 87170 3606
rect 85776 3466 86066 3482
rect 85764 3460 86066 3466
rect 85816 3454 86066 3460
rect 85764 3402 85816 3408
rect 86868 3324 86920 3330
rect 86868 3266 86920 3272
rect 86880 480 86908 3266
rect 74970 326 75408 354
rect 74970 -960 75082 326
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87800 218 87828 3674
rect 99012 3664 99064 3670
rect 96816 3602 97106 3618
rect 109408 3664 109460 3670
rect 99064 3612 99314 3618
rect 99012 3606 99314 3612
rect 109408 3606 109460 3612
rect 96804 3596 97106 3602
rect 96856 3590 97106 3596
rect 99024 3590 99314 3606
rect 102232 3596 102284 3602
rect 96804 3538 96856 3544
rect 102232 3538 102284 3544
rect 92388 3528 92440 3534
rect 92440 3476 92690 3482
rect 92388 3470 92690 3476
rect 90364 3460 90416 3466
rect 92400 3454 92690 3470
rect 90364 3402 90416 3408
rect 89536 3392 89588 3398
rect 89536 3334 89588 3340
rect 87984 3194 88274 3210
rect 87972 3188 88274 3194
rect 88024 3182 88274 3188
rect 87972 3130 88024 3136
rect 89076 3120 89128 3126
rect 89128 3068 89378 3074
rect 89076 3062 89378 3068
rect 89088 3046 89378 3062
rect 87942 218 88054 480
rect 87800 190 88054 218
rect 87942 -960 88054 190
rect 89138 354 89250 480
rect 89548 354 89576 3334
rect 90376 480 90404 3402
rect 96252 3392 96304 3398
rect 96252 3334 96304 3340
rect 93952 3256 94004 3262
rect 93952 3198 94004 3204
rect 90468 2990 90496 3060
rect 91296 3046 91586 3074
rect 93504 3058 93794 3074
rect 93492 3052 93794 3058
rect 90456 2984 90508 2990
rect 90456 2926 90508 2932
rect 91296 2854 91324 3046
rect 93544 3046 93794 3052
rect 93492 2994 93544 3000
rect 91560 2984 91612 2990
rect 91560 2926 91612 2932
rect 91284 2848 91336 2854
rect 91284 2790 91336 2796
rect 91572 480 91600 2926
rect 92756 2848 92808 2854
rect 92756 2790 92808 2796
rect 92768 480 92796 2790
rect 93964 480 93992 3198
rect 95148 3052 95200 3058
rect 95148 2994 95200 3000
rect 95160 480 95188 2994
rect 95988 2922 96016 3060
rect 95976 2916 96028 2922
rect 95976 2858 96028 2864
rect 96264 480 96292 3334
rect 100128 3330 100418 3346
rect 100116 3324 100418 3330
rect 100168 3318 100418 3324
rect 100116 3266 100168 3272
rect 101036 3188 101088 3194
rect 101036 3130 101088 3136
rect 98736 3120 98788 3126
rect 98736 3062 98788 3068
rect 97448 2916 97500 2922
rect 97448 2858 97500 2864
rect 97460 480 97488 2858
rect 98644 2848 98696 2854
rect 98644 2790 98696 2796
rect 98656 1290 98684 2790
rect 98644 1284 98696 1290
rect 98644 1226 98696 1232
rect 98748 1170 98776 3062
rect 99840 2848 99892 2854
rect 99840 2790 99892 2796
rect 98656 1142 98776 1170
rect 98656 480 98684 1142
rect 99852 480 99880 2790
rect 101048 480 101076 3130
rect 102244 480 102272 3538
rect 103612 3528 103664 3534
rect 102336 3466 102626 3482
rect 103664 3476 103730 3482
rect 103612 3470 103730 3476
rect 102324 3460 102626 3466
rect 102376 3454 102626 3460
rect 103624 3454 103730 3470
rect 105728 3460 105780 3466
rect 102324 3402 102376 3408
rect 105728 3402 105780 3408
rect 103336 3324 103388 3330
rect 103336 3266 103388 3272
rect 103348 480 103376 3266
rect 104544 3046 104834 3074
rect 104544 2990 104572 3046
rect 104532 2984 104584 2990
rect 104532 2926 104584 2932
rect 104624 2984 104676 2990
rect 104624 2926 104676 2932
rect 104636 1578 104664 2926
rect 104544 1550 104664 1578
rect 104544 480 104572 1550
rect 105740 480 105768 3402
rect 109040 3392 109092 3398
rect 109092 3340 109250 3346
rect 109040 3334 109250 3340
rect 109052 3318 109250 3334
rect 106740 3256 106792 3262
rect 107200 3256 107252 3262
rect 106792 3204 107042 3210
rect 106740 3198 107042 3204
rect 107200 3198 107252 3204
rect 106752 3182 107042 3198
rect 105924 1290 105952 3060
rect 107212 1714 107240 3198
rect 107856 3058 108146 3074
rect 107844 3052 108146 3058
rect 107896 3046 108146 3052
rect 108488 3052 108540 3058
rect 107844 2994 107896 3000
rect 108488 2994 108540 3000
rect 106936 1686 107240 1714
rect 105912 1284 105964 1290
rect 105912 1226 105964 1232
rect 106936 480 106964 1686
rect 89138 326 89576 354
rect 89138 -960 89250 326
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 354 108202 480
rect 108500 354 108528 2994
rect 109420 1850 109448 3606
rect 110512 3528 110564 3534
rect 110512 3470 110564 3476
rect 110064 3046 110354 3074
rect 110064 2922 110092 3046
rect 110052 2916 110104 2922
rect 110052 2858 110104 2864
rect 109328 1822 109448 1850
rect 109328 480 109356 1822
rect 110524 480 110552 3470
rect 112812 3392 112864 3398
rect 112812 3334 112864 3340
rect 111156 3120 111208 3126
rect 111616 3120 111668 3126
rect 111208 3068 111458 3074
rect 111156 3062 111458 3068
rect 111616 3062 111668 3068
rect 111168 3046 111458 3062
rect 111628 480 111656 3062
rect 112548 2854 112576 3060
rect 112536 2848 112588 2854
rect 112536 2790 112588 2796
rect 112824 480 112852 3334
rect 113100 3194 113666 3210
rect 113088 3188 113666 3194
rect 113140 3182 113666 3188
rect 113088 3130 113140 3136
rect 114020 480 114048 3742
rect 116400 3732 116452 3738
rect 116400 3674 116452 3680
rect 114480 3602 114770 3618
rect 114468 3596 114770 3602
rect 114520 3590 114770 3596
rect 114468 3538 114520 3544
rect 115584 3330 115874 3346
rect 115572 3324 115874 3330
rect 115624 3318 115874 3324
rect 115572 3266 115624 3272
rect 115204 2916 115256 2922
rect 115204 2858 115256 2864
rect 115216 480 115244 2858
rect 116412 480 116440 3674
rect 121184 3664 121236 3670
rect 121236 3612 121394 3618
rect 121184 3606 121394 3612
rect 121092 3596 121144 3602
rect 121196 3590 121394 3606
rect 121092 3538 121144 3544
rect 117792 3466 118082 3482
rect 117780 3460 118082 3466
rect 117832 3454 118082 3460
rect 117780 3402 117832 3408
rect 117596 3324 117648 3330
rect 117596 3266 117648 3272
rect 116964 2990 116992 3060
rect 116952 2984 117004 2990
rect 116952 2926 117004 2932
rect 117608 480 117636 3266
rect 118608 3256 118660 3262
rect 119896 3256 119948 3262
rect 118660 3204 119186 3210
rect 118608 3198 119186 3204
rect 119896 3198 119948 3204
rect 118620 3182 119186 3198
rect 118792 2848 118844 2854
rect 118792 2790 118844 2796
rect 118804 480 118832 2790
rect 119908 480 119936 3198
rect 120000 3058 120290 3074
rect 119988 3052 120290 3058
rect 120040 3046 120290 3052
rect 119988 2994 120040 3000
rect 121104 480 121132 3538
rect 122300 480 122328 3810
rect 125508 3800 125560 3806
rect 125560 3748 125810 3754
rect 125508 3742 125810 3748
rect 125520 3726 125810 3742
rect 127728 3738 128018 3754
rect 127716 3732 128018 3738
rect 127768 3726 128018 3732
rect 127716 3674 127768 3680
rect 125048 3664 125100 3670
rect 135444 3664 135496 3670
rect 125048 3606 125100 3612
rect 122380 3528 122432 3534
rect 122432 3476 122498 3482
rect 122380 3470 122498 3476
rect 122392 3454 122498 3470
rect 124128 3392 124180 3398
rect 124180 3340 124706 3346
rect 124128 3334 124706 3340
rect 124140 3318 124706 3334
rect 123300 3120 123352 3126
rect 123352 3068 123602 3074
rect 123300 3062 123602 3068
rect 123312 3046 123602 3062
rect 123484 2984 123536 2990
rect 123484 2926 123536 2932
rect 123496 480 123524 2926
rect 108090 326 108528 354
rect 108090 -960 108202 326
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 354 124762 480
rect 125060 354 125088 3606
rect 132144 3602 132434 3618
rect 143632 3664 143684 3670
rect 135496 3612 135746 3618
rect 135444 3606 135746 3612
rect 153108 3664 153160 3670
rect 143632 3606 143684 3612
rect 132132 3596 132434 3602
rect 132184 3590 132434 3596
rect 135456 3590 135746 3606
rect 136456 3596 136508 3602
rect 132132 3538 132184 3544
rect 136456 3538 136508 3544
rect 127072 3528 127124 3534
rect 127072 3470 127124 3476
rect 125968 3392 126020 3398
rect 125968 3334 126020 3340
rect 125980 1714 126008 3334
rect 126900 2922 126928 3060
rect 126888 2916 126940 2922
rect 126888 2858 126940 2864
rect 127084 1850 127112 3470
rect 131764 3460 131816 3466
rect 131764 3402 131816 3408
rect 128832 3330 129122 3346
rect 128820 3324 129122 3330
rect 128872 3318 129122 3324
rect 129372 3324 129424 3330
rect 128820 3266 128872 3272
rect 129372 3266 129424 3272
rect 128176 3052 128228 3058
rect 128176 2994 128228 3000
rect 125888 1686 126008 1714
rect 126992 1822 127112 1850
rect 125888 480 125916 1686
rect 126992 480 127020 1822
rect 128188 480 128216 2994
rect 129384 480 129412 3266
rect 131028 3256 131080 3262
rect 131080 3204 131330 3210
rect 131028 3198 131330 3204
rect 131040 3182 131330 3198
rect 130212 2854 130240 3060
rect 130568 2984 130620 2990
rect 130568 2926 130620 2932
rect 130200 2848 130252 2854
rect 130200 2790 130252 2796
rect 130580 480 130608 2926
rect 131776 480 131804 3402
rect 134352 3194 134642 3210
rect 134340 3188 134642 3194
rect 134392 3182 134642 3188
rect 134340 3130 134392 3136
rect 134156 3120 134208 3126
rect 134156 3062 134208 3068
rect 132960 2916 133012 2922
rect 132960 2858 133012 2864
rect 132972 480 133000 2858
rect 134168 480 134196 3062
rect 135260 2848 135312 2854
rect 135260 2790 135312 2796
rect 135272 480 135300 2790
rect 136468 480 136496 3538
rect 137652 3528 137704 3534
rect 139216 3528 139268 3534
rect 137704 3476 137954 3482
rect 137652 3470 137954 3476
rect 139216 3470 139268 3476
rect 137664 3454 137954 3470
rect 136640 3392 136692 3398
rect 136692 3340 136850 3346
rect 136640 3334 136850 3340
rect 136652 3318 136850 3334
rect 137652 3188 137704 3194
rect 137652 3130 137704 3136
rect 137664 480 137692 3130
rect 138768 3058 139058 3074
rect 138756 3052 139058 3058
rect 138808 3046 139058 3052
rect 138756 2994 138808 3000
rect 124650 326 125088 354
rect 124650 -960 124762 326
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 354 138930 480
rect 139228 354 139256 3470
rect 142264 3466 142370 3482
rect 142252 3460 142370 3466
rect 142304 3454 142370 3460
rect 142528 3460 142580 3466
rect 142252 3402 142304 3408
rect 142528 3402 142580 3408
rect 139872 3330 140162 3346
rect 139860 3324 140162 3330
rect 139912 3318 140162 3324
rect 139860 3266 139912 3272
rect 140044 3256 140096 3262
rect 140044 3198 140096 3204
rect 140056 480 140084 3198
rect 140976 3046 141266 3074
rect 140976 2990 141004 3046
rect 140964 2984 141016 2990
rect 140964 2926 141016 2932
rect 141240 2984 141292 2990
rect 141240 2926 141292 2932
rect 141252 480 141280 2926
rect 142540 1578 142568 3402
rect 143184 3058 143474 3074
rect 143172 3052 143474 3058
rect 143224 3046 143474 3052
rect 143172 2994 143224 3000
rect 143644 1850 143672 3606
rect 146496 3602 146786 3618
rect 153160 3612 153410 3618
rect 153108 3606 153410 3612
rect 146484 3596 146786 3602
rect 146536 3590 146786 3596
rect 149520 3596 149572 3602
rect 146484 3538 146536 3544
rect 153120 3590 153410 3606
rect 158640 3602 158930 3618
rect 158628 3596 158930 3602
rect 149520 3538 149572 3544
rect 158680 3590 158930 3596
rect 158628 3538 158680 3544
rect 148692 3528 148744 3534
rect 148744 3476 148994 3482
rect 148692 3470 148994 3476
rect 148704 3454 148994 3470
rect 148324 3324 148376 3330
rect 148324 3266 148376 3272
rect 147784 3194 147890 3210
rect 147772 3188 147890 3194
rect 147824 3182 147890 3188
rect 147772 3130 147824 3136
rect 144276 3120 144328 3126
rect 147128 3120 147180 3126
rect 144328 3068 144578 3074
rect 144276 3062 144578 3068
rect 144288 3046 144578 3062
rect 145392 3046 145682 3074
rect 147128 3062 147180 3068
rect 145932 3052 145984 3058
rect 144736 2916 144788 2922
rect 144736 2858 144788 2864
rect 142448 1550 142568 1578
rect 143552 1822 143672 1850
rect 142448 480 142476 1550
rect 143552 480 143580 1822
rect 144748 480 144776 2858
rect 145392 2854 145420 3046
rect 145932 2994 145984 3000
rect 145380 2848 145432 2854
rect 145380 2790 145432 2796
rect 145944 480 145972 2994
rect 147140 480 147168 3062
rect 148336 480 148364 3266
rect 149532 480 149560 3538
rect 153016 3528 153068 3534
rect 151740 3466 152306 3482
rect 153016 3470 153068 3476
rect 160192 3528 160244 3534
rect 160192 3470 160244 3476
rect 151728 3460 152306 3466
rect 151780 3454 152306 3460
rect 151728 3402 151780 3408
rect 149796 3392 149848 3398
rect 149848 3340 150098 3346
rect 149796 3334 150098 3340
rect 149808 3318 150098 3334
rect 150912 3046 151202 3074
rect 151820 3052 151872 3058
rect 150912 2990 150940 3046
rect 151820 2994 151872 3000
rect 150900 2984 150952 2990
rect 150900 2926 150952 2932
rect 150624 2916 150676 2922
rect 150624 2858 150676 2864
rect 150636 480 150664 2858
rect 151832 480 151860 2994
rect 153028 480 153056 3470
rect 155776 3460 155828 3466
rect 155776 3402 155828 3408
rect 154028 3256 154080 3262
rect 154028 3198 154080 3204
rect 138818 326 139256 354
rect 138818 -960 138930 326
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154040 218 154068 3198
rect 155316 3120 155368 3126
rect 154224 3046 154514 3074
rect 155368 3068 155618 3074
rect 155316 3062 155618 3068
rect 155328 3046 155618 3062
rect 154224 2854 154252 3046
rect 154212 2848 154264 2854
rect 154212 2790 154264 2796
rect 154182 218 154294 480
rect 154040 190 154294 218
rect 154182 -960 154294 190
rect 155378 354 155490 480
rect 155788 354 155816 3402
rect 157260 3330 157826 3346
rect 157248 3324 157826 3330
rect 157300 3318 157826 3324
rect 158168 3324 158220 3330
rect 157248 3266 157300 3272
rect 158168 3266 158220 3272
rect 156432 3194 156722 3210
rect 156420 3188 156722 3194
rect 156472 3182 156722 3188
rect 156420 3130 156472 3136
rect 156604 2984 156656 2990
rect 156604 2926 156656 2932
rect 156616 480 156644 2926
rect 155378 326 155816 354
rect 155378 -960 155490 326
rect 156574 -960 156686 480
rect 157770 354 157882 480
rect 158180 354 158208 3266
rect 160204 3262 160232 3470
rect 166080 3460 166132 3466
rect 166080 3402 166132 3408
rect 161296 3324 161348 3330
rect 161296 3266 161348 3272
rect 160192 3256 160244 3262
rect 160192 3198 160244 3204
rect 160020 2922 160048 3060
rect 160848 3058 161138 3074
rect 160836 3052 161138 3058
rect 160888 3046 161138 3052
rect 160836 2994 160888 3000
rect 160008 2916 160060 2922
rect 160008 2858 160060 2864
rect 160100 2916 160152 2922
rect 160100 2858 160152 2864
rect 158904 2848 158956 2854
rect 158904 2790 158956 2796
rect 158916 480 158944 2790
rect 160112 480 160140 2858
rect 161308 480 161336 3266
rect 161940 3256 161992 3262
rect 163688 3256 163740 3262
rect 161992 3204 162242 3210
rect 161940 3198 162242 3204
rect 163688 3198 163740 3204
rect 161952 3182 162242 3198
rect 162768 3120 162820 3126
rect 162820 3068 163346 3074
rect 162768 3062 163346 3068
rect 162492 3052 162544 3058
rect 162780 3046 163346 3062
rect 162492 2994 162544 3000
rect 162504 480 162532 2994
rect 163700 480 163728 3198
rect 164160 3194 164450 3210
rect 164148 3188 164450 3194
rect 164200 3182 164450 3188
rect 164148 3130 164200 3136
rect 164884 3120 164936 3126
rect 164884 3062 164936 3068
rect 164896 480 164924 3062
rect 165540 2990 165568 3060
rect 165528 2984 165580 2990
rect 165528 2926 165580 2932
rect 166092 480 166120 3402
rect 166356 3392 166408 3398
rect 174084 3392 174136 3398
rect 166408 3340 166658 3346
rect 166356 3334 166658 3340
rect 166368 3318 166658 3334
rect 169680 3330 169970 3346
rect 174136 3340 174386 3346
rect 174084 3334 174386 3340
rect 169668 3324 169970 3330
rect 169720 3318 169970 3324
rect 174096 3318 174386 3334
rect 181824 3330 182114 3346
rect 181812 3324 182114 3330
rect 169668 3266 169720 3272
rect 181864 3318 182114 3324
rect 564190 3330 564388 3346
rect 564190 3324 564400 3330
rect 564190 3318 564348 3324
rect 181812 3266 181864 3272
rect 564348 3266 564400 3272
rect 583392 3324 583444 3330
rect 583392 3266 583444 3272
rect 171876 3256 171928 3262
rect 174268 3256 174320 3262
rect 171928 3204 172178 3210
rect 171876 3198 172178 3204
rect 180892 3256 180944 3262
rect 174268 3198 174320 3204
rect 170772 3188 170824 3194
rect 171888 3182 172178 3198
rect 170772 3130 170824 3136
rect 167184 2984 167236 2990
rect 167184 2926 167236 2932
rect 167196 480 167224 2926
rect 167748 2854 167776 3060
rect 168852 2922 168880 3060
rect 168840 2916 168892 2922
rect 168840 2858 168892 2864
rect 169576 2916 169628 2922
rect 169576 2858 169628 2864
rect 167736 2848 167788 2854
rect 167736 2790 167788 2796
rect 168380 2848 168432 2854
rect 168380 2790 168432 2796
rect 168392 480 168420 2790
rect 169588 480 169616 2858
rect 170784 480 170812 3130
rect 172980 3120 173032 3126
rect 170876 3058 171074 3074
rect 173440 3120 173492 3126
rect 173032 3068 173282 3074
rect 172980 3062 173282 3068
rect 173440 3062 173492 3068
rect 170864 3052 171074 3058
rect 170916 3046 171074 3052
rect 171968 3052 172020 3058
rect 170864 2994 170916 3000
rect 172992 3046 173282 3062
rect 171968 2994 172020 3000
rect 171980 480 172008 2994
rect 173452 1714 173480 3062
rect 173176 1686 173480 1714
rect 173176 480 173204 1686
rect 174280 480 174308 3198
rect 178512 3194 178802 3210
rect 184940 3256 184992 3262
rect 180944 3204 181010 3210
rect 180892 3198 181010 3204
rect 200304 3256 200356 3262
rect 184940 3198 184992 3204
rect 178500 3188 178802 3194
rect 178552 3182 178802 3188
rect 180904 3182 181010 3198
rect 181444 3188 181496 3194
rect 178500 3130 178552 3136
rect 181444 3130 181496 3136
rect 179052 3120 179104 3126
rect 175476 2990 175504 3060
rect 176304 3046 176594 3074
rect 179052 3062 179104 3068
rect 175464 2984 175516 2990
rect 175464 2926 175516 2932
rect 175832 2984 175884 2990
rect 175832 2926 175884 2932
rect 157770 326 158208 354
rect 157770 -960 157882 326
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 354 175546 480
rect 175844 354 175872 2926
rect 176304 2854 176332 3046
rect 177684 2922 177712 3060
rect 177856 2984 177908 2990
rect 177856 2926 177908 2932
rect 177672 2916 177724 2922
rect 177672 2858 177724 2864
rect 176292 2848 176344 2854
rect 176292 2790 176344 2796
rect 176660 1352 176712 1358
rect 176660 1294 176712 1300
rect 176672 480 176700 1294
rect 177868 480 177896 2926
rect 179064 480 179092 3062
rect 179616 3058 179906 3074
rect 179604 3052 179906 3058
rect 179656 3046 179906 3052
rect 179604 2994 179656 3000
rect 180248 2848 180300 2854
rect 180248 2790 180300 2796
rect 180260 480 180288 2790
rect 181456 480 181484 3130
rect 182548 3052 182600 3058
rect 182548 2994 182600 3000
rect 182928 3046 183218 3074
rect 182560 480 182588 2994
rect 182928 2922 182956 3046
rect 182916 2916 182968 2922
rect 182916 2858 182968 2864
rect 183744 2916 183796 2922
rect 183744 2858 183796 2864
rect 183756 480 183784 2858
rect 184308 1358 184336 3060
rect 184296 1352 184348 1358
rect 184296 1294 184348 1300
rect 184952 480 184980 3198
rect 188448 3194 188738 3210
rect 188436 3188 188738 3194
rect 188488 3182 188738 3188
rect 189552 3182 189842 3210
rect 191760 3194 192050 3210
rect 206100 3256 206152 3262
rect 200304 3198 200356 3204
rect 191748 3188 192050 3194
rect 188436 3130 188488 3136
rect 186320 3120 186372 3126
rect 186372 3068 186530 3074
rect 186320 3062 186530 3068
rect 185412 2990 185440 3060
rect 186332 3046 186530 3062
rect 187344 3046 187634 3074
rect 189552 3058 189580 3182
rect 191800 3182 192050 3188
rect 195612 3188 195664 3194
rect 191748 3130 191800 3136
rect 195612 3130 195664 3136
rect 190552 3120 190604 3126
rect 190552 3062 190604 3068
rect 189540 3052 189592 3058
rect 185400 2984 185452 2990
rect 185400 2926 185452 2932
rect 187344 2854 187372 3046
rect 189540 2994 189592 3000
rect 189724 3052 189776 3058
rect 189724 2994 189776 3000
rect 187332 2848 187384 2854
rect 187332 2790 187384 2796
rect 187332 1352 187384 1358
rect 187332 1294 187384 1300
rect 186136 1216 186188 1222
rect 186136 1158 186188 1164
rect 186148 480 186176 1158
rect 187344 480 187372 1294
rect 188896 1284 188948 1290
rect 188896 1226 188948 1232
rect 175434 326 175872 354
rect 175434 -960 175546 326
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 354 188610 480
rect 188908 354 188936 1226
rect 189736 480 189764 2994
rect 188498 326 188936 354
rect 188498 -960 188610 326
rect 189694 -960 189806 480
rect 190564 354 190592 3062
rect 190656 3046 190946 3074
rect 190656 2922 190684 3046
rect 190644 2916 190696 2922
rect 190644 2858 190696 2864
rect 192392 2916 192444 2922
rect 192392 2858 192444 2864
rect 190798 354 190910 480
rect 190564 326 190910 354
rect 190798 -960 190910 326
rect 191994 354 192106 480
rect 192404 354 192432 2858
rect 193140 1222 193168 3060
rect 193220 2780 193272 2786
rect 193220 2722 193272 2728
rect 193128 1216 193180 1222
rect 193128 1158 193180 1164
rect 193232 480 193260 2722
rect 194244 1358 194272 3060
rect 194416 2984 194468 2990
rect 194416 2926 194468 2932
rect 194232 1352 194284 1358
rect 194232 1294 194284 1300
rect 194428 480 194456 2926
rect 195348 1290 195376 3060
rect 195336 1284 195388 1290
rect 195336 1226 195388 1232
rect 195624 480 195652 3130
rect 197268 3120 197320 3126
rect 196176 3058 196466 3074
rect 197320 3068 197570 3074
rect 197268 3062 197570 3068
rect 196164 3052 196466 3058
rect 196216 3046 196466 3052
rect 197280 3046 197570 3062
rect 198384 3046 198674 3074
rect 199488 3046 199778 3074
rect 196164 2994 196216 3000
rect 198384 2922 198412 3046
rect 199108 2984 199160 2990
rect 199108 2926 199160 2932
rect 198372 2916 198424 2922
rect 198372 2858 198424 2864
rect 198280 1352 198332 1358
rect 198280 1294 198332 1300
rect 197176 1284 197228 1290
rect 197176 1226 197228 1232
rect 191994 326 192432 354
rect 191994 -960 192106 326
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 354 196890 480
rect 197188 354 197216 1226
rect 196778 326 197216 354
rect 197882 354 197994 480
rect 198292 354 198320 1294
rect 199120 480 199148 2926
rect 199488 2854 199516 3046
rect 199476 2848 199528 2854
rect 199476 2790 199528 2796
rect 200316 480 200344 3198
rect 201696 3194 201986 3210
rect 556712 3256 556764 3262
rect 206152 3204 206402 3210
rect 206100 3198 206402 3204
rect 201684 3188 201986 3194
rect 201736 3182 201986 3188
rect 206112 3182 206402 3198
rect 224880 3194 225170 3210
rect 220268 3188 220320 3194
rect 201684 3130 201736 3136
rect 220268 3130 220320 3136
rect 224868 3188 225170 3194
rect 224920 3182 225170 3188
rect 556462 3204 556712 3210
rect 575112 3256 575164 3262
rect 556462 3198 556764 3204
rect 556462 3182 556752 3198
rect 560878 3194 561168 3210
rect 575112 3198 575164 3204
rect 560878 3188 561180 3194
rect 560878 3182 561128 3188
rect 224868 3130 224920 3136
rect 561128 3130 561180 3136
rect 202696 3120 202748 3126
rect 200592 3058 200882 3074
rect 208308 3120 208360 3126
rect 202696 3062 202748 3068
rect 200580 3052 200882 3058
rect 200632 3046 200882 3052
rect 200580 2994 200632 3000
rect 201500 2916 201552 2922
rect 201500 2858 201552 2864
rect 201512 480 201540 2858
rect 202708 480 202736 3062
rect 203076 1290 203104 3060
rect 203892 3052 203944 3058
rect 203892 2994 203944 3000
rect 203064 1284 203116 1290
rect 203064 1226 203116 1232
rect 203904 480 203932 2994
rect 204180 1358 204208 3060
rect 205008 3046 205298 3074
rect 206940 3046 207506 3074
rect 209872 3120 209924 3126
rect 208360 3068 208610 3074
rect 208308 3062 208610 3068
rect 208320 3046 208610 3062
rect 209424 3058 209714 3074
rect 214932 3120 214984 3126
rect 209872 3062 209924 3068
rect 209412 3052 209714 3058
rect 205008 2990 205036 3046
rect 206940 2990 206968 3046
rect 209464 3046 209714 3052
rect 209412 2994 209464 3000
rect 204996 2984 205048 2990
rect 204996 2926 205048 2932
rect 206928 2984 206980 2990
rect 206928 2926 206980 2932
rect 208584 2984 208636 2990
rect 208584 2926 208636 2932
rect 206192 2916 206244 2922
rect 206192 2858 206244 2864
rect 205088 2848 205140 2854
rect 205088 2790 205140 2796
rect 204168 1352 204220 1358
rect 204168 1294 204220 1300
rect 205100 480 205128 2790
rect 206204 480 206232 2858
rect 207388 1352 207440 1358
rect 207388 1294 207440 1300
rect 207400 480 207428 1294
rect 208596 480 208624 2926
rect 209884 1578 209912 3062
rect 210528 3046 210818 3074
rect 211632 3046 211922 3074
rect 212172 3052 212224 3058
rect 210528 2854 210556 3046
rect 211632 2922 211660 3046
rect 212172 2994 212224 3000
rect 211620 2916 211672 2922
rect 211620 2858 211672 2864
rect 210516 2848 210568 2854
rect 210516 2790 210568 2796
rect 210976 2848 211028 2854
rect 210976 2790 211028 2796
rect 209792 1550 209912 1578
rect 209792 480 209820 1550
rect 210988 480 211016 2790
rect 212184 480 212212 2994
rect 213012 1358 213040 3060
rect 213840 3046 214130 3074
rect 215668 3120 215720 3126
rect 214984 3068 215234 3074
rect 214932 3062 215234 3068
rect 215668 3062 215720 3068
rect 214944 3046 215234 3062
rect 213840 2990 213868 3046
rect 213828 2984 213880 2990
rect 213828 2926 213880 2932
rect 214472 2984 214524 2990
rect 214472 2926 214524 2932
rect 213368 2916 213420 2922
rect 213368 2858 213420 2864
rect 213000 1352 213052 1358
rect 213000 1294 213052 1300
rect 213380 480 213408 2858
rect 214484 480 214512 2926
rect 215680 480 215708 3062
rect 216048 3046 216338 3074
rect 217152 3058 217442 3074
rect 217140 3052 217442 3058
rect 216048 2854 216076 3046
rect 217192 3046 217442 3052
rect 217980 3046 218546 3074
rect 219256 3052 219308 3058
rect 217140 2994 217192 3000
rect 217980 2922 218008 3046
rect 219256 2994 219308 3000
rect 219360 3046 219650 3074
rect 217968 2916 218020 2922
rect 217968 2858 218020 2864
rect 218060 2916 218112 2922
rect 218060 2858 218112 2864
rect 216036 2848 216088 2854
rect 216036 2790 216088 2796
rect 216864 2848 216916 2854
rect 216864 2790 216916 2796
rect 216876 480 216904 2790
rect 218072 480 218100 2858
rect 219268 480 219296 2994
rect 219360 2990 219388 3046
rect 219348 2984 219400 2990
rect 219348 2926 219400 2932
rect 197882 326 198320 354
rect 196778 -960 196890 326
rect 197882 -960 197994 326
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220280 218 220308 3130
rect 220452 3120 220504 3126
rect 221556 3120 221608 3126
rect 220504 3068 220754 3074
rect 220452 3062 220754 3068
rect 225972 3120 226024 3126
rect 221556 3062 221608 3068
rect 220464 3046 220754 3062
rect 221568 480 221596 3062
rect 221844 2854 221872 3060
rect 222948 2922 222976 3060
rect 223500 3058 224066 3074
rect 228732 3120 228784 3126
rect 226024 3068 226274 3074
rect 225972 3062 226274 3068
rect 223488 3052 224066 3058
rect 223540 3046 224066 3052
rect 225984 3046 226274 3062
rect 223488 2994 223540 3000
rect 223948 2984 224000 2990
rect 223948 2926 224000 2932
rect 225144 2984 225196 2990
rect 225144 2926 225196 2932
rect 222936 2916 222988 2922
rect 222936 2858 222988 2864
rect 223120 2916 223172 2922
rect 223120 2858 223172 2864
rect 221832 2848 221884 2854
rect 221832 2790 221884 2796
rect 220422 218 220534 480
rect 220280 190 220534 218
rect 220422 -960 220534 190
rect 221526 -960 221638 480
rect 222722 354 222834 480
rect 223132 354 223160 2858
rect 223960 480 223988 2926
rect 225156 480 225184 2926
rect 227364 2922 227392 3060
rect 228192 3058 228482 3074
rect 228732 3062 228784 3068
rect 232596 3120 232648 3126
rect 239312 3120 239364 3126
rect 232648 3068 232898 3074
rect 232596 3062 232898 3068
rect 228180 3052 228482 3058
rect 228232 3046 228482 3052
rect 228180 2994 228232 3000
rect 227352 2916 227404 2922
rect 227352 2858 227404 2864
rect 227536 2916 227588 2922
rect 227536 2858 227588 2864
rect 226340 2848 226392 2854
rect 226340 2790 226392 2796
rect 226352 480 226380 2790
rect 227548 480 227576 2858
rect 228744 480 228772 3062
rect 229572 2990 229600 3060
rect 229836 3052 229888 3058
rect 229836 2994 229888 3000
rect 229560 2984 229612 2990
rect 229560 2926 229612 2932
rect 229848 480 229876 2994
rect 230676 2854 230704 3060
rect 231032 2984 231084 2990
rect 231032 2926 231084 2932
rect 230664 2848 230716 2854
rect 230664 2790 230716 2796
rect 231044 480 231072 2926
rect 231780 2922 231808 3060
rect 232608 3046 232898 3062
rect 233712 3058 234002 3074
rect 233700 3052 234002 3058
rect 233752 3046 234002 3052
rect 234620 3052 234672 3058
rect 233700 2994 233752 3000
rect 234620 2994 234672 3000
rect 231768 2916 231820 2922
rect 231768 2858 231820 2864
rect 232228 2916 232280 2922
rect 232228 2858 232280 2864
rect 232240 480 232268 2858
rect 233424 2848 233476 2854
rect 233424 2790 233476 2796
rect 233436 480 233464 2790
rect 234632 480 234660 2994
rect 235092 2990 235120 3060
rect 235080 2984 235132 2990
rect 235080 2926 235132 2932
rect 235816 2984 235868 2990
rect 235816 2926 235868 2932
rect 235828 480 235856 2926
rect 236196 2922 236224 3060
rect 236184 2916 236236 2922
rect 236184 2858 236236 2864
rect 237012 2916 237064 2922
rect 237012 2858 237064 2864
rect 237024 480 237052 2858
rect 237300 2854 237328 3060
rect 238128 3058 238418 3074
rect 239312 3062 239364 3068
rect 242532 3120 242584 3126
rect 543464 3120 543516 3126
rect 242584 3068 242834 3074
rect 242532 3062 242834 3068
rect 238116 3052 238418 3058
rect 238168 3046 238418 3052
rect 238116 2994 238168 3000
rect 237288 2848 237340 2854
rect 237288 2790 237340 2796
rect 238116 2848 238168 2854
rect 238116 2790 238168 2796
rect 238128 480 238156 2790
rect 239324 480 239352 3062
rect 239508 2990 239536 3060
rect 240508 3052 240560 3058
rect 240508 2994 240560 3000
rect 239496 2984 239548 2990
rect 239496 2926 239548 2932
rect 240520 480 240548 2994
rect 240612 2922 240640 3060
rect 240600 2916 240652 2922
rect 240600 2858 240652 2864
rect 241716 2854 241744 3060
rect 242544 3046 242834 3062
rect 243648 3058 243938 3074
rect 243636 3052 243938 3058
rect 243688 3046 243938 3052
rect 243636 2994 243688 3000
rect 245028 2990 245056 3060
rect 245200 3052 245252 3058
rect 245200 2994 245252 3000
rect 242072 2984 242124 2990
rect 242072 2926 242124 2932
rect 245016 2984 245068 2990
rect 245016 2926 245068 2932
rect 241704 2848 241756 2854
rect 241704 2790 241756 2796
rect 222722 326 223160 354
rect 222722 -960 222834 326
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 354 241786 480
rect 242084 354 242112 2926
rect 244096 2916 244148 2922
rect 244096 2858 244148 2864
rect 242900 2848 242952 2854
rect 242900 2790 242952 2796
rect 242912 480 242940 2790
rect 244108 480 244136 2858
rect 245212 480 245240 2994
rect 246132 2854 246160 3060
rect 247236 2922 247264 3060
rect 248064 3058 248354 3074
rect 248052 3052 248354 3058
rect 248104 3046 248354 3052
rect 248788 3052 248840 3058
rect 248052 2994 248104 3000
rect 248788 2994 248840 3000
rect 247592 2984 247644 2990
rect 247592 2926 247644 2932
rect 247224 2916 247276 2922
rect 247224 2858 247276 2864
rect 246120 2848 246172 2854
rect 246120 2790 246172 2796
rect 246396 2848 246448 2854
rect 246396 2790 246448 2796
rect 246408 480 246436 2790
rect 247604 480 247632 2926
rect 248800 480 248828 2994
rect 249444 2854 249472 3060
rect 250548 2990 250576 3060
rect 251376 3058 251666 3074
rect 251364 3052 251666 3058
rect 251416 3046 251666 3052
rect 251364 2994 251416 3000
rect 250536 2984 250588 2990
rect 250536 2926 250588 2932
rect 252756 2922 252784 3060
rect 253480 2984 253532 2990
rect 253480 2926 253532 2932
rect 249984 2916 250036 2922
rect 249984 2858 250036 2864
rect 252744 2916 252796 2922
rect 252744 2858 252796 2864
rect 249432 2848 249484 2854
rect 249432 2790 249484 2796
rect 249996 480 250024 2858
rect 252376 2848 252428 2854
rect 252376 2790 252428 2796
rect 251180 808 251232 814
rect 251180 750 251232 756
rect 251192 480 251220 750
rect 252388 480 252416 2790
rect 253492 480 253520 2926
rect 253860 814 253888 3060
rect 254676 2916 254728 2922
rect 254676 2858 254728 2864
rect 253848 808 253900 814
rect 253848 750 253900 756
rect 254688 480 254716 2858
rect 254964 2854 254992 3060
rect 256068 2990 256096 3060
rect 256056 2984 256108 2990
rect 256056 2926 256108 2932
rect 257172 2922 257200 3060
rect 257160 2916 257212 2922
rect 257160 2858 257212 2864
rect 258276 2854 258304 3060
rect 254952 2848 255004 2854
rect 254952 2790 255004 2796
rect 255872 2848 255924 2854
rect 255872 2790 255924 2796
rect 258264 2848 258316 2854
rect 258264 2790 258316 2796
rect 255884 480 255912 2790
rect 259380 1358 259408 3060
rect 257068 1352 257120 1358
rect 257068 1294 257120 1300
rect 259368 1352 259420 1358
rect 259368 1294 259420 1300
rect 259460 1352 259512 1358
rect 259460 1294 259512 1300
rect 257080 480 257108 1294
rect 258264 1284 258316 1290
rect 258264 1226 258316 1232
rect 258276 480 258304 1226
rect 259472 480 259500 1294
rect 260484 1290 260512 3060
rect 260656 2848 260708 2854
rect 260656 2790 260708 2796
rect 260472 1284 260524 1290
rect 260472 1226 260524 1232
rect 260668 480 260696 2790
rect 261588 1358 261616 3060
rect 261760 2916 261812 2922
rect 261760 2858 261812 2864
rect 261576 1352 261628 1358
rect 261576 1294 261628 1300
rect 261772 480 261800 2858
rect 262692 2854 262720 3060
rect 263796 2922 263824 3060
rect 263784 2916 263836 2922
rect 263784 2858 263836 2864
rect 262680 2848 262732 2854
rect 262680 2790 262732 2796
rect 264900 1358 264928 3060
rect 262956 1352 263008 1358
rect 262956 1294 263008 1300
rect 264888 1352 264940 1358
rect 264888 1294 264940 1300
rect 265348 1352 265400 1358
rect 265348 1294 265400 1300
rect 262968 480 262996 1294
rect 264152 1284 264204 1290
rect 264152 1226 264204 1232
rect 264164 480 264192 1226
rect 265360 480 265388 1294
rect 266004 1290 266032 3060
rect 267108 1358 267136 3060
rect 267096 1352 267148 1358
rect 267096 1294 267148 1300
rect 267740 1352 267792 1358
rect 267740 1294 267792 1300
rect 265992 1284 266044 1290
rect 265992 1226 266044 1232
rect 266544 1284 266596 1290
rect 266544 1226 266596 1232
rect 266556 480 266584 1226
rect 267752 480 267780 1294
rect 268212 1290 268240 3060
rect 269316 1358 269344 3060
rect 269304 1352 269356 1358
rect 269304 1294 269356 1300
rect 268200 1284 268252 1290
rect 268200 1226 268252 1232
rect 270040 1284 270092 1290
rect 270040 1226 270092 1232
rect 268844 1216 268896 1222
rect 268844 1158 268896 1164
rect 268856 480 268884 1158
rect 270052 480 270080 1226
rect 270420 1222 270448 3060
rect 271236 1352 271288 1358
rect 271236 1294 271288 1300
rect 270408 1216 270460 1222
rect 270408 1158 270460 1164
rect 271248 480 271276 1294
rect 271524 1290 271552 3060
rect 272628 1358 272656 3060
rect 272616 1352 272668 1358
rect 272616 1294 272668 1300
rect 273628 1352 273680 1358
rect 273628 1294 273680 1300
rect 271512 1284 271564 1290
rect 271512 1226 271564 1232
rect 272432 1284 272484 1290
rect 272432 1226 272484 1232
rect 272444 480 272472 1226
rect 273640 480 273668 1294
rect 273732 1290 273760 3060
rect 274836 1358 274864 3060
rect 275296 3046 275954 3074
rect 276124 3046 277058 3074
rect 274824 1352 274876 1358
rect 274824 1294 274876 1300
rect 273720 1284 273772 1290
rect 273720 1226 273772 1232
rect 241674 326 242112 354
rect 241674 -960 241786 326
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 354 274906 480
rect 275296 354 275324 3046
rect 276124 1578 276152 3046
rect 276032 1550 276152 1578
rect 276032 480 276060 1550
rect 278148 1358 278176 3060
rect 278792 3046 279266 3074
rect 277124 1352 277176 1358
rect 277124 1294 277176 1300
rect 278136 1352 278188 1358
rect 278136 1294 278188 1300
rect 277136 480 277164 1294
rect 274794 326 275324 354
rect 274794 -960 274906 326
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 354 278402 480
rect 278792 354 278820 3046
rect 280356 1358 280384 3060
rect 281184 3046 281474 3074
rect 281920 3046 282578 3074
rect 283392 3046 283682 3074
rect 284312 3046 284786 3074
rect 285416 3046 285890 3074
rect 279516 1352 279568 1358
rect 279516 1294 279568 1300
rect 280344 1352 280396 1358
rect 280344 1294 280396 1300
rect 279528 480 279556 1294
rect 278290 326 278820 354
rect 278290 -960 278402 326
rect 279486 -960 279598 480
rect 280682 354 280794 480
rect 281184 354 281212 3046
rect 281920 480 281948 3046
rect 280682 326 281212 354
rect 280682 -960 280794 326
rect 281878 -960 281990 480
rect 283074 354 283186 480
rect 283392 354 283420 3046
rect 284312 480 284340 3046
rect 285416 480 285444 3046
rect 283074 326 283420 354
rect 283074 -960 283186 326
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 354 286682 480
rect 286980 354 287008 3060
rect 287808 3046 288098 3074
rect 287808 480 287836 3046
rect 286570 326 287008 354
rect 286570 -960 286682 326
rect 287766 -960 287878 480
rect 288962 354 289074 480
rect 289188 354 289216 3060
rect 290200 3046 290306 3074
rect 290200 480 290228 3046
rect 291396 480 291424 3060
rect 292592 480 292620 3060
rect 293696 480 293724 3060
rect 294814 3046 294920 3074
rect 295918 3046 296116 3074
rect 297022 3046 297312 3074
rect 294892 480 294920 3046
rect 296088 480 296116 3046
rect 297284 480 297312 3046
rect 288962 326 289216 354
rect 288962 -960 289074 326
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298112 354 298140 3060
rect 299230 3046 299704 3074
rect 300334 3046 300808 3074
rect 301438 3046 301728 3074
rect 302542 3046 303200 3074
rect 303646 3046 303936 3074
rect 299676 480 299704 3046
rect 300780 480 300808 3046
rect 298438 354 298550 480
rect 298112 326 298550 354
rect 298438 -960 298550 326
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301700 354 301728 3046
rect 303172 480 303200 3046
rect 301934 354 302046 480
rect 301700 326 302046 354
rect 301934 -960 302046 326
rect 303130 -960 303242 480
rect 303908 354 303936 3046
rect 304736 2854 304764 3060
rect 305854 3046 306328 3074
rect 304724 2848 304776 2854
rect 304724 2790 304776 2796
rect 305552 2848 305604 2854
rect 305552 2790 305604 2796
rect 305564 480 305592 2790
rect 304326 354 304438 480
rect 303908 326 304438 354
rect 304326 -960 304438 326
rect 305522 -960 305634 480
rect 306300 354 306328 3046
rect 306944 2854 306972 3060
rect 308062 3046 308996 3074
rect 306932 2848 306984 2854
rect 306932 2790 306984 2796
rect 307944 2848 307996 2854
rect 307944 2790 307996 2796
rect 307956 480 307984 2790
rect 308968 1578 308996 3046
rect 309152 2854 309180 3060
rect 310256 2990 310284 3060
rect 310244 2984 310296 2990
rect 310244 2926 310296 2932
rect 311360 2854 311388 3060
rect 311440 2984 311492 2990
rect 311440 2926 311492 2932
rect 309140 2848 309192 2854
rect 309140 2790 309192 2796
rect 310244 2848 310296 2854
rect 310244 2790 310296 2796
rect 311348 2848 311400 2854
rect 311348 2790 311400 2796
rect 308968 1550 309088 1578
rect 309060 480 309088 1550
rect 310256 480 310284 2790
rect 311452 480 311480 2926
rect 312464 2922 312492 3060
rect 312452 2916 312504 2922
rect 312452 2858 312504 2864
rect 313568 2854 313596 3060
rect 314580 2922 314608 3060
rect 313832 2916 313884 2922
rect 313832 2858 313884 2864
rect 314568 2916 314620 2922
rect 314568 2858 314620 2864
rect 312636 2848 312688 2854
rect 312636 2790 312688 2796
rect 313556 2848 313608 2854
rect 313556 2790 313608 2796
rect 312648 480 312676 2790
rect 313844 480 313872 2858
rect 315776 2854 315804 3060
rect 316880 2922 316908 3060
rect 316224 2916 316276 2922
rect 316224 2858 316276 2864
rect 316868 2916 316920 2922
rect 316868 2858 316920 2864
rect 315028 2848 315080 2854
rect 315028 2790 315080 2796
rect 315764 2848 315816 2854
rect 315764 2790 315816 2796
rect 315040 480 315068 2790
rect 316236 480 316264 2858
rect 317984 2854 318012 3060
rect 319088 2922 319116 3060
rect 318524 2916 318576 2922
rect 318524 2858 318576 2864
rect 319076 2916 319128 2922
rect 319076 2858 319128 2864
rect 317328 2848 317380 2854
rect 317328 2790 317380 2796
rect 317972 2848 318024 2854
rect 317972 2790 318024 2796
rect 317340 480 317368 2790
rect 318536 480 318564 2858
rect 320100 2854 320128 3060
rect 321296 2922 321324 3060
rect 320916 2916 320968 2922
rect 320916 2858 320968 2864
rect 321284 2916 321336 2922
rect 321284 2858 321336 2864
rect 319720 2848 319772 2854
rect 319720 2790 319772 2796
rect 320088 2848 320140 2854
rect 320088 2790 320140 2796
rect 319732 480 319760 2790
rect 320928 480 320956 2858
rect 322400 2854 322428 3060
rect 323504 2922 323532 3060
rect 323308 2916 323360 2922
rect 323308 2858 323360 2864
rect 323492 2916 323544 2922
rect 323492 2858 323544 2864
rect 322112 2848 322164 2854
rect 322112 2790 322164 2796
rect 322388 2848 322440 2854
rect 322388 2790 322440 2796
rect 322124 480 322152 2790
rect 323320 480 323348 2858
rect 324608 2854 324636 3060
rect 325712 2990 325740 3060
rect 326830 3046 327028 3074
rect 325700 2984 325752 2990
rect 325700 2926 325752 2932
rect 325608 2916 325660 2922
rect 325608 2858 325660 2864
rect 324412 2848 324464 2854
rect 324412 2790 324464 2796
rect 324596 2848 324648 2854
rect 324596 2790 324648 2796
rect 324424 480 324452 2790
rect 325620 480 325648 2858
rect 327000 2854 327028 3046
rect 327920 2922 327948 3060
rect 329024 2990 329052 3060
rect 328000 2984 328052 2990
rect 328000 2926 328052 2932
rect 329012 2984 329064 2990
rect 329012 2926 329064 2932
rect 327908 2916 327960 2922
rect 327908 2858 327960 2864
rect 326804 2848 326856 2854
rect 326804 2790 326856 2796
rect 326988 2848 327040 2854
rect 326988 2790 327040 2796
rect 326816 480 326844 2790
rect 328012 480 328040 2926
rect 330128 2854 330156 3060
rect 331140 2922 331168 3060
rect 332336 2990 332364 3060
rect 333454 3058 333744 3074
rect 333454 3052 333756 3058
rect 333454 3046 333704 3052
rect 333704 2994 333756 3000
rect 331588 2984 331640 2990
rect 331588 2926 331640 2932
rect 332324 2984 332376 2990
rect 332324 2926 332376 2932
rect 330392 2916 330444 2922
rect 330392 2858 330444 2864
rect 331128 2916 331180 2922
rect 331128 2858 331180 2864
rect 329196 2848 329248 2854
rect 329196 2790 329248 2796
rect 330116 2848 330168 2854
rect 330116 2790 330168 2796
rect 329208 480 329236 2790
rect 330404 480 330432 2858
rect 331600 480 331628 2926
rect 334544 2922 334572 3060
rect 335084 2984 335136 2990
rect 335084 2926 335136 2932
rect 333888 2916 333940 2922
rect 333888 2858 333940 2864
rect 334532 2916 334584 2922
rect 334532 2858 334584 2864
rect 332692 2848 332744 2854
rect 332692 2790 332744 2796
rect 332704 480 332732 2790
rect 333900 480 333928 2858
rect 335096 480 335124 2926
rect 335648 2854 335676 3060
rect 336280 3052 336332 3058
rect 336280 2994 336332 3000
rect 335636 2848 335688 2854
rect 335636 2790 335688 2796
rect 336292 480 336320 2994
rect 336660 1358 336688 3060
rect 337476 2916 337528 2922
rect 337476 2858 337528 2864
rect 336648 1352 336700 1358
rect 336648 1294 336700 1300
rect 337488 480 337516 2858
rect 337856 882 337884 3060
rect 338960 2854 338988 3060
rect 340064 2922 340092 3060
rect 341168 2990 341196 3060
rect 341156 2984 341208 2990
rect 341156 2926 341208 2932
rect 340052 2916 340104 2922
rect 340052 2858 340104 2864
rect 338672 2848 338724 2854
rect 338672 2790 338724 2796
rect 338948 2848 339000 2854
rect 338948 2790 339000 2796
rect 342076 2848 342128 2854
rect 342076 2790 342128 2796
rect 337844 876 337896 882
rect 337844 818 337896 824
rect 338684 480 338712 2790
rect 339868 1352 339920 1358
rect 339868 1294 339920 1300
rect 339880 480 339908 1294
rect 342088 1170 342116 2790
rect 342180 1358 342208 3060
rect 342996 2916 343048 2922
rect 342996 2858 343048 2864
rect 342168 1352 342220 1358
rect 342168 1294 342220 1300
rect 342088 1142 342208 1170
rect 340972 876 341024 882
rect 340972 818 341024 824
rect 340984 480 341012 818
rect 342180 480 342208 1142
rect 306718 354 306830 480
rect 306300 326 306830 354
rect 306718 -960 306830 326
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343008 354 343036 2858
rect 343376 1290 343404 3060
rect 344494 3046 344784 3074
rect 344560 2984 344612 2990
rect 344560 2926 344612 2932
rect 343364 1284 343416 1290
rect 343364 1226 343416 1232
rect 344572 480 344600 2926
rect 343334 354 343446 480
rect 343008 326 343446 354
rect 343334 -960 343446 326
rect 344530 -960 344642 480
rect 344756 66 344784 3046
rect 345584 1018 345612 3060
rect 346688 2854 346716 3060
rect 346676 2848 346728 2854
rect 346676 2790 346728 2796
rect 345756 1352 345808 1358
rect 345756 1294 345808 1300
rect 345572 1012 345624 1018
rect 345572 954 345624 960
rect 345768 480 345796 1294
rect 346952 1284 347004 1290
rect 346952 1226 347004 1232
rect 346964 480 346992 1226
rect 347700 882 347728 3060
rect 348896 1358 348924 3060
rect 348884 1352 348936 1358
rect 348884 1294 348936 1300
rect 350000 1290 350028 3060
rect 350448 2848 350500 2854
rect 350448 2790 350500 2796
rect 349988 1284 350040 1290
rect 349988 1226 350040 1232
rect 349252 1012 349304 1018
rect 349252 954 349304 960
rect 347688 876 347740 882
rect 347688 818 347740 824
rect 349264 480 349292 954
rect 350460 480 350488 2790
rect 351104 1018 351132 3060
rect 352208 1154 352236 3060
rect 353220 2854 353248 3060
rect 353208 2848 353260 2854
rect 353208 2790 353260 2796
rect 352840 1352 352892 1358
rect 352840 1294 352892 1300
rect 352196 1148 352248 1154
rect 352196 1090 352248 1096
rect 351092 1012 351144 1018
rect 351092 954 351144 960
rect 351644 876 351696 882
rect 351644 818 351696 824
rect 351656 480 351684 818
rect 352852 480 352880 1294
rect 354036 1284 354088 1290
rect 354036 1226 354088 1232
rect 354048 480 354076 1226
rect 344744 60 344796 66
rect 344744 2 344796 8
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 82 348138 480
rect 348026 66 348280 82
rect 348026 60 348292 66
rect 348026 54 348240 60
rect 348026 -960 348138 54
rect 348240 2 348292 8
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 354416 270 354444 3060
rect 355520 1086 355548 3060
rect 356624 1358 356652 3060
rect 357532 2848 357584 2854
rect 357532 2790 357584 2796
rect 356612 1352 356664 1358
rect 356612 1294 356664 1300
rect 356336 1148 356388 1154
rect 356336 1090 356388 1096
rect 355508 1080 355560 1086
rect 355508 1022 355560 1028
rect 355232 1012 355284 1018
rect 355232 954 355284 960
rect 355244 480 355272 954
rect 356348 480 356376 1090
rect 357544 480 357572 2790
rect 357728 1290 357756 3060
rect 357716 1284 357768 1290
rect 357716 1226 357768 1232
rect 358740 950 358768 3060
rect 359936 1222 359964 3060
rect 359924 1216 359976 1222
rect 359924 1158 359976 1164
rect 361040 1154 361068 3060
rect 361120 1352 361172 1358
rect 361120 1294 361172 1300
rect 361028 1148 361080 1154
rect 361028 1090 361080 1096
rect 359924 1080 359976 1086
rect 359924 1022 359976 1028
rect 358728 944 358780 950
rect 358728 886 358780 892
rect 359936 480 359964 1022
rect 361132 480 361160 1294
rect 362144 1018 362172 3060
rect 362316 1284 362368 1290
rect 362316 1226 362368 1232
rect 362132 1012 362184 1018
rect 362132 954 362184 960
rect 362328 480 362356 1226
rect 354404 264 354456 270
rect 354404 206 354456 212
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 218 358810 480
rect 358912 264 358964 270
rect 358698 212 358912 218
rect 358698 206 358964 212
rect 358698 190 358952 206
rect 358698 -960 358810 190
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363248 66 363276 3060
rect 364260 1358 364288 3060
rect 364248 1352 364300 1358
rect 364248 1294 364300 1300
rect 365456 1290 365484 3060
rect 365444 1284 365496 1290
rect 365444 1226 365496 1232
rect 366560 1222 366588 3060
rect 364616 1216 364668 1222
rect 364616 1158 364668 1164
rect 366548 1216 366600 1222
rect 366548 1158 366600 1164
rect 363512 944 363564 950
rect 363512 886 363564 892
rect 363524 480 363552 886
rect 364628 480 364656 1158
rect 367664 1154 367692 3060
rect 365444 1148 365496 1154
rect 365444 1090 365496 1096
rect 367652 1148 367704 1154
rect 367652 1090 367704 1096
rect 363236 60 363288 66
rect 363236 2 363288 8
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365456 354 365484 1090
rect 367008 1012 367060 1018
rect 367008 954 367060 960
rect 367020 480 367048 954
rect 368768 882 368796 3060
rect 369400 1352 369452 1358
rect 369400 1294 369452 1300
rect 368756 876 368808 882
rect 368756 818 368808 824
rect 369412 480 369440 1294
rect 369780 1018 369808 3060
rect 370976 1290 371004 3060
rect 372094 3046 372384 3074
rect 372356 2854 372384 3046
rect 372344 2848 372396 2854
rect 372344 2790 372396 2796
rect 370228 1284 370280 1290
rect 370228 1226 370280 1232
rect 370964 1284 371016 1290
rect 370964 1226 371016 1232
rect 369768 1012 369820 1018
rect 369768 954 369820 960
rect 365782 354 365894 480
rect 365456 326 365894 354
rect 365782 -960 365894 326
rect 366978 -960 367090 480
rect 368174 82 368286 480
rect 367848 66 368286 82
rect 367836 60 368286 66
rect 367888 54 368286 60
rect 367836 2 367888 8
rect 368174 -960 368286 54
rect 369370 -960 369482 480
rect 370240 354 370268 1226
rect 371332 1216 371384 1222
rect 371332 1158 371384 1164
rect 370566 354 370678 480
rect 370240 326 370678 354
rect 371344 354 371372 1158
rect 372896 1148 372948 1154
rect 372896 1090 372948 1096
rect 372908 480 372936 1090
rect 373184 1086 373212 3060
rect 374288 1358 374316 3060
rect 374276 1352 374328 1358
rect 374276 1294 374328 1300
rect 375300 1154 375328 3060
rect 376116 1284 376168 1290
rect 376116 1226 376168 1232
rect 375288 1148 375340 1154
rect 375288 1090 375340 1096
rect 373172 1080 373224 1086
rect 373172 1022 373224 1028
rect 375288 1012 375340 1018
rect 375288 954 375340 960
rect 373908 876 373960 882
rect 373908 818 373960 824
rect 371670 354 371782 480
rect 371344 326 371782 354
rect 370566 -960 370678 326
rect 371670 -960 371782 326
rect 372866 -960 372978 480
rect 373920 354 373948 818
rect 375300 480 375328 954
rect 374062 354 374174 480
rect 373920 326 374174 354
rect 374062 -960 374174 326
rect 375258 -960 375370 480
rect 376128 354 376156 1226
rect 376496 1018 376524 3060
rect 377600 1290 377628 3060
rect 377680 2848 377732 2854
rect 377680 2790 377732 2796
rect 377588 1284 377640 1290
rect 377588 1226 377640 1232
rect 376484 1012 376536 1018
rect 376484 954 376536 960
rect 377692 480 377720 2790
rect 378704 1222 378732 3060
rect 379612 1352 379664 1358
rect 379612 1294 379664 1300
rect 378692 1216 378744 1222
rect 378692 1158 378744 1164
rect 378508 1080 378560 1086
rect 378508 1022 378560 1028
rect 376454 354 376566 480
rect 376128 326 376566 354
rect 376454 -960 376566 326
rect 377650 -960 377762 480
rect 378520 354 378548 1022
rect 378846 354 378958 480
rect 378520 326 378958 354
rect 379624 354 379652 1294
rect 379808 1154 379836 3060
rect 379796 1148 379848 1154
rect 379796 1090 379848 1096
rect 379950 354 380062 480
rect 379624 326 380062 354
rect 378846 -960 378958 326
rect 379950 -960 380062 326
rect 380820 270 380848 3060
rect 381176 1080 381228 1086
rect 381176 1022 381228 1028
rect 381188 480 381216 1022
rect 380808 264 380860 270
rect 380808 206 380860 212
rect 381146 -960 381258 480
rect 382016 474 382044 3060
rect 382372 1012 382424 1018
rect 382372 954 382424 960
rect 382384 480 382412 954
rect 382004 468 382056 474
rect 382004 410 382056 416
rect 382342 -960 382454 480
rect 383120 66 383148 3060
rect 384224 1358 384252 3060
rect 384212 1352 384264 1358
rect 384212 1294 384264 1300
rect 383568 1284 383620 1290
rect 383568 1226 383620 1232
rect 383580 480 383608 1226
rect 384396 1216 384448 1222
rect 384396 1158 384448 1164
rect 383108 60 383160 66
rect 383108 2 383160 8
rect 383538 -960 383650 480
rect 384408 354 384436 1158
rect 385328 1086 385356 3060
rect 386340 1154 386368 3060
rect 387536 1222 387564 3060
rect 388640 1290 388668 3060
rect 388628 1284 388680 1290
rect 388628 1226 388680 1232
rect 387524 1216 387576 1222
rect 387524 1158 387576 1164
rect 385960 1148 386012 1154
rect 385960 1090 386012 1096
rect 386328 1148 386380 1154
rect 386328 1090 386380 1096
rect 385316 1080 385368 1086
rect 385316 1022 385368 1028
rect 385972 480 386000 1090
rect 389744 610 389772 3060
rect 390652 1352 390704 1358
rect 390652 1294 390704 1300
rect 389732 604 389784 610
rect 389732 546 389784 552
rect 390664 480 390692 1294
rect 384734 354 384846 480
rect 384408 326 384846 354
rect 384734 -960 384846 326
rect 385930 -960 386042 480
rect 386788 264 386840 270
rect 387126 218 387238 480
rect 387892 468 387944 474
rect 387892 410 387944 416
rect 387904 354 387932 410
rect 388230 354 388342 480
rect 387904 326 388342 354
rect 386840 212 387238 218
rect 386788 206 387238 212
rect 386800 190 387238 206
rect 387126 -960 387238 190
rect 388230 -960 388342 326
rect 389426 82 389538 480
rect 389426 66 389680 82
rect 389426 60 389692 66
rect 389426 54 389640 60
rect 389426 -960 389538 54
rect 389640 2 389692 8
rect 390622 -960 390734 480
rect 390848 66 390876 3060
rect 391676 3046 391874 3074
rect 391676 270 391704 3046
rect 392676 1148 392728 1154
rect 392676 1090 392728 1096
rect 391848 1080 391900 1086
rect 391848 1022 391900 1028
rect 391860 480 391888 1022
rect 391664 264 391716 270
rect 391664 206 391716 212
rect 390836 60 390888 66
rect 390836 2 390888 8
rect 391818 -960 391930 480
rect 392688 354 392716 1090
rect 393056 678 393084 3060
rect 394160 1086 394188 3060
rect 395264 1222 395292 3060
rect 396368 1358 396396 3060
rect 396356 1352 396408 1358
rect 396356 1294 396408 1300
rect 395344 1284 395396 1290
rect 395344 1226 395396 1232
rect 394240 1216 394292 1222
rect 394240 1158 394292 1164
rect 395252 1216 395304 1222
rect 395252 1158 395304 1164
rect 394148 1080 394200 1086
rect 394148 1022 394200 1028
rect 393044 672 393096 678
rect 393044 614 393096 620
rect 394252 480 394280 1158
rect 395356 480 395384 1226
rect 397380 1154 397408 3060
rect 397368 1148 397420 1154
rect 397368 1090 397420 1096
rect 396540 604 396592 610
rect 396540 546 396592 552
rect 396552 480 396580 546
rect 393014 354 393126 480
rect 392688 326 393126 354
rect 393014 -960 393126 326
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 82 397818 480
rect 398576 338 398604 3060
rect 398564 332 398616 338
rect 398564 274 398616 280
rect 398748 264 398800 270
rect 398902 218 399014 480
rect 398800 212 399014 218
rect 398748 206 399014 212
rect 398760 190 399014 206
rect 397706 66 397960 82
rect 397706 60 397972 66
rect 397706 54 397920 60
rect 397706 -960 397818 54
rect 397920 2 397972 8
rect 398902 -960 399014 190
rect 399680 134 399708 3060
rect 400784 678 400812 3060
rect 401324 1080 401376 1086
rect 401324 1022 401376 1028
rect 400128 672 400180 678
rect 400128 614 400180 620
rect 400772 672 400824 678
rect 400772 614 400824 620
rect 400140 480 400168 614
rect 401336 480 401364 1022
rect 401888 746 401916 3060
rect 402520 1216 402572 1222
rect 402520 1158 402572 1164
rect 401876 740 401928 746
rect 401876 682 401928 688
rect 402532 480 402560 1158
rect 399668 128 399720 134
rect 399668 70 399720 76
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 402900 66 402928 3060
rect 403624 1352 403676 1358
rect 403624 1294 403676 1300
rect 403636 480 403664 1294
rect 404096 1290 404124 3060
rect 404084 1284 404136 1290
rect 404084 1226 404136 1232
rect 404820 1148 404872 1154
rect 404820 1090 404872 1096
rect 404832 480 404860 1090
rect 402888 60 402940 66
rect 402888 2 402940 8
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405200 270 405228 3060
rect 406304 1358 406332 3060
rect 406292 1352 406344 1358
rect 406292 1294 406344 1300
rect 405986 354 406098 480
rect 405986 338 406240 354
rect 405986 332 406252 338
rect 405986 326 406200 332
rect 405188 264 405240 270
rect 405188 206 405240 212
rect 405986 -960 406098 326
rect 406200 274 406252 280
rect 407028 128 407080 134
rect 407182 82 407294 480
rect 407408 406 407436 3060
rect 408420 610 408448 3060
rect 409236 740 409288 746
rect 409236 682 409288 688
rect 408592 672 408644 678
rect 408592 614 408644 620
rect 408408 604 408460 610
rect 408408 546 408460 552
rect 407396 400 407448 406
rect 407396 342 407448 348
rect 407080 76 407294 82
rect 407028 70 407294 76
rect 407040 54 407294 70
rect 407182 -960 407294 54
rect 408378 218 408490 480
rect 408604 218 408632 614
rect 408378 190 408632 218
rect 409248 218 409276 682
rect 409616 678 409644 3060
rect 410734 3046 411024 3074
rect 411838 3046 412128 3074
rect 409604 672 409656 678
rect 409604 614 409656 620
rect 409574 218 409686 480
rect 409248 190 409686 218
rect 408378 -960 408490 190
rect 409574 -960 409686 190
rect 410770 82 410882 480
rect 410996 338 411024 3046
rect 411904 1284 411956 1290
rect 411904 1226 411956 1232
rect 411916 480 411944 1226
rect 410984 332 411036 338
rect 410984 274 411036 280
rect 410770 66 411024 82
rect 410770 60 411036 66
rect 410770 54 410984 60
rect 410770 -960 410882 54
rect 410984 2 411036 8
rect 411874 -960 411986 480
rect 412100 474 412128 3046
rect 412928 1222 412956 3060
rect 413940 1290 413968 3060
rect 414296 1352 414348 1358
rect 414296 1294 414348 1300
rect 413928 1284 413980 1290
rect 413928 1226 413980 1232
rect 412916 1216 412968 1222
rect 412916 1158 412968 1164
rect 414308 480 414336 1294
rect 415136 1086 415164 3060
rect 415124 1080 415176 1086
rect 415124 1022 415176 1028
rect 416240 950 416268 3060
rect 416228 944 416280 950
rect 416228 886 416280 892
rect 416688 604 416740 610
rect 416688 546 416740 552
rect 416700 480 416728 546
rect 412088 468 412140 474
rect 412088 410 412140 416
rect 412824 264 412876 270
rect 413070 218 413182 480
rect 412876 212 413182 218
rect 412824 206 413182 212
rect 412836 190 413182 206
rect 413070 -960 413182 190
rect 414266 -960 414378 480
rect 415308 400 415360 406
rect 415462 354 415574 480
rect 415360 348 415574 354
rect 415308 342 415574 348
rect 415320 326 415574 342
rect 415462 -960 415574 326
rect 416658 -960 416770 480
rect 417344 66 417372 3060
rect 417884 672 417936 678
rect 417884 614 417936 620
rect 417896 480 417924 614
rect 417332 60 417384 66
rect 417332 2 417384 8
rect 417854 -960 417966 480
rect 418448 202 418476 3060
rect 419460 1358 419488 3060
rect 419448 1352 419500 1358
rect 419448 1294 419500 1300
rect 420656 1154 420684 3060
rect 421760 1222 421788 3060
rect 422576 1284 422628 1290
rect 422576 1226 422628 1232
rect 421380 1216 421432 1222
rect 421380 1158 421432 1164
rect 421748 1216 421800 1222
rect 421748 1158 421800 1164
rect 420644 1148 420696 1154
rect 420644 1090 420696 1096
rect 421392 480 421420 1158
rect 422588 480 422616 1226
rect 422864 1018 422892 3060
rect 423404 1080 423456 1086
rect 423404 1022 423456 1028
rect 422852 1012 422904 1018
rect 422852 954 422904 960
rect 418958 354 419070 480
rect 418632 338 419070 354
rect 418620 332 419070 338
rect 418672 326 419070 332
rect 418620 274 418672 280
rect 418436 196 418488 202
rect 418436 138 418488 144
rect 418958 -960 419070 326
rect 420154 354 420266 480
rect 420368 468 420420 474
rect 420368 410 420420 416
rect 420380 354 420408 410
rect 420154 326 420408 354
rect 420154 -960 420266 326
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423416 354 423444 1022
rect 423742 354 423854 480
rect 423416 326 423854 354
rect 423742 -960 423854 326
rect 423968 134 423996 3060
rect 424980 1086 425008 3060
rect 426176 1290 426204 3060
rect 426164 1284 426216 1290
rect 426164 1226 426216 1232
rect 424968 1080 425020 1086
rect 424968 1022 425020 1028
rect 424968 944 425020 950
rect 424968 886 425020 892
rect 424980 480 425008 886
rect 427280 814 427308 3060
rect 428384 1358 428412 3060
rect 428280 1352 428332 1358
rect 428280 1294 428332 1300
rect 428372 1352 428424 1358
rect 428372 1294 428424 1300
rect 427268 808 427320 814
rect 427268 750 427320 756
rect 428292 762 428320 1294
rect 429292 1148 429344 1154
rect 429292 1090 429344 1096
rect 428292 734 428504 762
rect 428476 480 428504 734
rect 423956 128 424008 134
rect 423956 70 424008 76
rect 424938 -960 425050 480
rect 426134 82 426246 480
rect 427238 218 427350 480
rect 426912 202 427350 218
rect 426900 196 427350 202
rect 426952 190 427350 196
rect 426900 138 426952 144
rect 425808 66 426246 82
rect 425796 60 426246 66
rect 425848 54 426246 60
rect 425796 2 425848 8
rect 426134 -960 426246 54
rect 427238 -960 427350 190
rect 428434 -960 428546 480
rect 429304 354 429332 1090
rect 429488 746 429516 3060
rect 429476 740 429528 746
rect 429476 682 429528 688
rect 430500 542 430528 3060
rect 430856 1216 430908 1222
rect 430856 1158 430908 1164
rect 430488 536 430540 542
rect 429630 354 429742 480
rect 430488 478 430540 484
rect 430868 480 430896 1158
rect 431696 610 431724 3060
rect 432800 1018 432828 3060
rect 431868 1012 431920 1018
rect 431868 954 431920 960
rect 432788 1012 432840 1018
rect 432788 954 432840 960
rect 431684 604 431736 610
rect 431684 546 431736 552
rect 429304 326 429742 354
rect 429630 -960 429742 326
rect 430826 -960 430938 480
rect 431880 354 431908 954
rect 433904 950 433932 3060
rect 435008 1154 435036 3060
rect 436020 1358 436048 3060
rect 436008 1352 436060 1358
rect 436008 1294 436060 1300
rect 435180 1284 435232 1290
rect 435180 1226 435232 1232
rect 434996 1148 435048 1154
rect 434996 1090 435048 1096
rect 434076 1080 434128 1086
rect 434076 1022 434128 1028
rect 433892 944 433944 950
rect 433892 886 433944 892
rect 432022 354 432134 480
rect 431880 326 432134 354
rect 432022 -960 432134 326
rect 433218 82 433330 480
rect 434088 354 434116 1022
rect 434414 354 434526 480
rect 434088 326 434526 354
rect 435192 354 435220 1226
rect 436744 808 436796 814
rect 436744 750 436796 756
rect 436756 480 436784 750
rect 435518 354 435630 480
rect 435192 326 435630 354
rect 433432 128 433484 134
rect 433218 76 433432 82
rect 433218 70 433484 76
rect 433218 54 433472 70
rect 433218 -960 433330 54
rect 434414 -960 434526 326
rect 435518 -960 435630 326
rect 436714 -960 436826 480
rect 437216 474 437244 3060
rect 438320 1290 438348 3060
rect 437572 1284 437624 1290
rect 437572 1226 437624 1232
rect 438308 1284 438360 1290
rect 438308 1226 438360 1232
rect 437204 468 437256 474
rect 437204 410 437256 416
rect 437584 354 437612 1226
rect 439424 1222 439452 3060
rect 439412 1216 439464 1222
rect 439412 1158 439464 1164
rect 440528 746 440556 3060
rect 441540 1086 441568 3060
rect 441528 1080 441580 1086
rect 441528 1022 441580 1028
rect 442632 1012 442684 1018
rect 442632 954 442684 960
rect 439136 740 439188 746
rect 439136 682 439188 688
rect 440516 740 440568 746
rect 440516 682 440568 688
rect 439148 480 439176 682
rect 441528 672 441580 678
rect 441528 614 441580 620
rect 440332 604 440384 610
rect 440332 546 440384 552
rect 440344 480 440372 546
rect 441540 480 441568 614
rect 442644 480 442672 954
rect 442736 814 442764 3060
rect 443840 1358 443868 3060
rect 444958 3046 445248 3074
rect 443828 1352 443880 1358
rect 443828 1294 443880 1300
rect 443552 1216 443604 1222
rect 443552 1158 443604 1164
rect 443564 1018 443592 1158
rect 445220 1154 445248 3046
rect 445852 1284 445904 1290
rect 445852 1226 445904 1232
rect 445024 1148 445076 1154
rect 445024 1090 445076 1096
rect 445208 1148 445260 1154
rect 445208 1090 445260 1096
rect 443552 1012 443604 1018
rect 443552 954 443604 960
rect 443460 944 443512 950
rect 443460 886 443512 892
rect 442724 808 442776 814
rect 442724 750 442776 756
rect 437910 354 438022 480
rect 437584 326 438022 354
rect 437910 -960 438022 326
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443472 354 443500 886
rect 445036 480 445064 1090
rect 443798 354 443910 480
rect 443472 326 443910 354
rect 443798 -960 443910 326
rect 444994 -960 445106 480
rect 445864 354 445892 1226
rect 446048 950 446076 3060
rect 446036 944 446088 950
rect 446036 886 446088 892
rect 447060 610 447088 3060
rect 448256 882 448284 3060
rect 449360 1290 449388 3060
rect 449348 1284 449400 1290
rect 449348 1226 449400 1232
rect 450464 1222 450492 3060
rect 448612 1216 448664 1222
rect 448612 1158 448664 1164
rect 450452 1216 450504 1222
rect 450452 1158 450504 1164
rect 448244 876 448296 882
rect 448244 818 448296 824
rect 447048 604 447100 610
rect 447048 546 447100 552
rect 447244 598 447456 626
rect 446190 354 446302 480
rect 447244 474 447272 598
rect 447428 480 447456 598
rect 448624 480 448652 1158
rect 449808 1012 449860 1018
rect 449808 954 449860 960
rect 449820 480 449848 954
rect 451568 746 451596 3060
rect 451740 1080 451792 1086
rect 451740 1022 451792 1028
rect 450912 740 450964 746
rect 450912 682 450964 688
rect 451556 740 451608 746
rect 451556 682 451608 688
rect 450924 480 450952 682
rect 447232 468 447284 474
rect 447232 410 447284 416
rect 445864 326 446302 354
rect 446190 -960 446302 326
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 451752 354 451780 1022
rect 452078 354 452190 480
rect 451752 326 452190 354
rect 452078 -960 452190 326
rect 452580 134 452608 3060
rect 453304 808 453356 814
rect 453304 750 453356 756
rect 453316 480 453344 750
rect 452568 128 452620 134
rect 452568 70 452620 76
rect 453274 -960 453386 480
rect 453776 338 453804 3060
rect 454132 1352 454184 1358
rect 454132 1294 454184 1300
rect 454144 354 454172 1294
rect 454880 1290 454908 3060
rect 454868 1284 454920 1290
rect 454868 1226 454920 1232
rect 455696 1148 455748 1154
rect 455696 1090 455748 1096
rect 455708 480 455736 1090
rect 455984 1086 456012 3060
rect 457088 1358 457116 3060
rect 457916 3046 458114 3074
rect 459310 3046 459508 3074
rect 460414 3046 460612 3074
rect 456984 1352 457036 1358
rect 456984 1294 457036 1300
rect 457076 1352 457128 1358
rect 457076 1294 457128 1300
rect 455972 1080 456024 1086
rect 455972 1022 456024 1028
rect 456892 944 456944 950
rect 456892 886 456944 892
rect 456904 480 456932 886
rect 456996 678 457024 1294
rect 456984 672 457036 678
rect 456984 614 457036 620
rect 454470 354 454582 480
rect 453764 332 453816 338
rect 454144 326 454582 354
rect 453764 274 453816 280
rect 454470 -960 454582 326
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 457916 270 457944 3046
rect 459192 876 459244 882
rect 459192 818 459244 824
rect 458088 604 458140 610
rect 458088 546 458140 552
rect 458100 480 458128 546
rect 459204 480 459232 818
rect 459480 542 459508 3046
rect 460020 672 460072 678
rect 460020 614 460072 620
rect 459468 536 459520 542
rect 457904 264 457956 270
rect 457904 206 457956 212
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 459468 478 459520 484
rect 460032 354 460060 614
rect 460358 354 460470 480
rect 460584 406 460612 3046
rect 461504 610 461532 3060
rect 462608 1290 462636 3060
rect 462596 1284 462648 1290
rect 462596 1226 462648 1232
rect 461584 1148 461636 1154
rect 461584 1090 461636 1096
rect 461492 604 461544 610
rect 461492 546 461544 552
rect 461596 480 461624 1090
rect 462412 808 462464 814
rect 462412 750 462464 756
rect 460032 326 460470 354
rect 460572 400 460624 406
rect 460572 342 460624 348
rect 460358 -960 460470 326
rect 461554 -960 461666 480
rect 462424 354 462452 750
rect 462750 354 462862 480
rect 462424 326 462862 354
rect 462750 -960 462862 326
rect 463620 66 463648 3060
rect 464816 678 464844 3060
rect 464804 672 464856 678
rect 464804 614 464856 620
rect 463946 82 464058 480
rect 465142 354 465254 480
rect 465000 338 465254 354
rect 464988 332 465254 338
rect 465040 326 465254 332
rect 464988 274 465040 280
rect 464160 128 464212 134
rect 463946 76 464160 82
rect 463946 70 464212 76
rect 463608 60 463660 66
rect 463608 2 463660 8
rect 463946 54 464200 70
rect 463946 -960 464058 54
rect 465142 -960 465254 326
rect 465828 202 465856 3060
rect 465908 1216 465960 1222
rect 465908 1158 465960 1164
rect 465920 354 465948 1158
rect 466246 354 466358 480
rect 465920 326 466358 354
rect 465816 196 465868 202
rect 465816 138 465868 144
rect 466246 -960 466358 326
rect 467024 134 467052 3060
rect 467472 1080 467524 1086
rect 467472 1022 467524 1028
rect 467484 480 467512 1022
rect 468128 746 468156 3060
rect 468300 1352 468352 1358
rect 468300 1294 468352 1300
rect 468116 740 468168 746
rect 468116 682 468168 688
rect 467012 128 467064 134
rect 467012 70 467064 76
rect 467442 -960 467554 480
rect 468312 354 468340 1294
rect 469140 1154 469168 3060
rect 469128 1148 469180 1154
rect 469128 1090 469180 1096
rect 468638 354 468750 480
rect 468312 326 468750 354
rect 468638 -960 468750 326
rect 469834 218 469946 480
rect 470336 474 470364 3060
rect 470784 536 470836 542
rect 470784 478 470836 484
rect 470324 468 470376 474
rect 470324 410 470376 416
rect 470796 354 470824 478
rect 471030 354 471142 480
rect 470796 326 471142 354
rect 471440 338 471468 3060
rect 472226 354 472338 480
rect 472440 400 472492 406
rect 472226 348 472440 354
rect 472226 342 472492 348
rect 470048 264 470100 270
rect 469834 212 470048 218
rect 469834 206 470100 212
rect 469834 190 470088 206
rect 469834 -960 469946 190
rect 471030 -960 471142 326
rect 471428 332 471480 338
rect 471428 274 471480 280
rect 472226 326 472480 342
rect 472226 -960 472338 326
rect 472544 270 472572 3060
rect 473452 604 473504 610
rect 473452 546 473504 552
rect 473464 480 473492 546
rect 473648 542 473676 3060
rect 474188 1284 474240 1290
rect 474188 1226 474240 1232
rect 473636 536 473688 542
rect 472532 264 472584 270
rect 472532 206 472584 212
rect 473422 -960 473534 480
rect 473636 478 473688 484
rect 474200 354 474228 1226
rect 474660 1086 474688 3060
rect 475856 1222 475884 3060
rect 476974 3046 477264 3074
rect 478078 3046 478368 3074
rect 475844 1216 475896 1222
rect 475844 1158 475896 1164
rect 474648 1080 474700 1086
rect 474648 1022 474700 1028
rect 476948 672 477000 678
rect 476948 614 477000 620
rect 476960 480 476988 614
rect 474526 354 474638 480
rect 474200 326 474638 354
rect 474526 -960 474638 326
rect 475722 82 475834 480
rect 475722 66 475976 82
rect 475722 60 475988 66
rect 475722 54 475936 60
rect 475722 -960 475834 54
rect 475936 2 475988 8
rect 476918 -960 477030 480
rect 477236 66 477264 3046
rect 478114 218 478226 480
rect 478340 406 478368 3046
rect 478328 400 478380 406
rect 478328 342 478380 348
rect 478114 202 478368 218
rect 479168 202 479196 3060
rect 480180 1290 480208 3060
rect 481376 1358 481404 3060
rect 481364 1352 481416 1358
rect 481364 1294 481416 1300
rect 480168 1284 480220 1290
rect 480168 1226 480220 1232
rect 481364 1148 481416 1154
rect 481364 1090 481416 1096
rect 480536 740 480588 746
rect 480536 682 480588 688
rect 480548 480 480576 682
rect 478114 196 478380 202
rect 478114 190 478328 196
rect 477224 60 477276 66
rect 477224 2 477276 8
rect 478114 -960 478226 190
rect 478328 138 478380 144
rect 479156 196 479208 202
rect 479156 138 479208 144
rect 478972 128 479024 134
rect 479310 82 479422 480
rect 479024 76 479422 82
rect 478972 70 479422 76
rect 478984 54 479422 70
rect 479310 -960 479422 54
rect 480506 -960 480618 480
rect 481376 354 481404 1090
rect 482480 746 482508 3060
rect 483584 814 483612 3060
rect 483572 808 483624 814
rect 483572 750 483624 756
rect 482468 740 482520 746
rect 482468 682 482520 688
rect 481702 354 481814 480
rect 482468 468 482520 474
rect 482468 410 482520 416
rect 481376 326 481814 354
rect 482480 354 482508 410
rect 482806 354 482918 480
rect 482480 326 482918 354
rect 481702 -960 481814 326
rect 482806 -960 482918 326
rect 484002 354 484114 480
rect 484688 474 484716 3060
rect 485700 882 485728 3060
rect 485688 876 485740 882
rect 485688 818 485740 824
rect 486896 678 486924 3060
rect 488000 1154 488028 3060
rect 488816 1216 488868 1222
rect 488816 1158 488868 1164
rect 487988 1148 488040 1154
rect 487988 1090 488040 1096
rect 487252 1080 487304 1086
rect 487252 1022 487304 1028
rect 486884 672 486936 678
rect 486884 614 486936 620
rect 486424 604 486476 610
rect 486424 546 486476 552
rect 486436 480 486464 546
rect 484676 468 484728 474
rect 484676 410 484728 416
rect 484002 338 484256 354
rect 484002 332 484268 338
rect 484002 326 484216 332
rect 484002 -960 484114 326
rect 484216 274 484268 280
rect 484860 264 484912 270
rect 485198 218 485310 480
rect 484912 212 485310 218
rect 484860 206 485310 212
rect 484872 190 485310 206
rect 485198 -960 485310 190
rect 486394 -960 486506 480
rect 487264 354 487292 1022
rect 488828 480 488856 1158
rect 489104 1018 489132 3060
rect 489092 1012 489144 1018
rect 489092 954 489144 960
rect 487590 354 487702 480
rect 487264 326 487702 354
rect 487590 -960 487702 326
rect 488786 -960 488898 480
rect 489890 82 490002 480
rect 490208 474 490236 3060
rect 491220 626 491248 3060
rect 492430 3046 492628 3074
rect 491220 598 491340 626
rect 490196 468 490248 474
rect 490196 410 490248 416
rect 490748 400 490800 406
rect 491086 354 491198 480
rect 490800 348 491198 354
rect 490748 342 491198 348
rect 490760 326 491198 342
rect 489890 66 490144 82
rect 489890 60 490156 66
rect 489890 54 490104 60
rect 489890 -960 490002 54
rect 490104 2 490156 8
rect 491086 -960 491198 326
rect 491312 134 491340 598
rect 492282 218 492394 480
rect 492282 202 492536 218
rect 492600 202 492628 3046
rect 493520 1290 493548 3060
rect 493140 1284 493192 1290
rect 493140 1226 493192 1232
rect 493508 1284 493560 1290
rect 493508 1226 493560 1232
rect 493152 354 493180 1226
rect 494624 950 494652 3060
rect 495728 1358 495756 3060
rect 494704 1352 494756 1358
rect 494704 1294 494756 1300
rect 495716 1352 495768 1358
rect 495716 1294 495768 1300
rect 494612 944 494664 950
rect 494612 886 494664 892
rect 494716 480 494744 1294
rect 495532 740 495584 746
rect 495532 682 495584 688
rect 493478 354 493590 480
rect 493152 326 493590 354
rect 492282 196 492548 202
rect 492282 190 492496 196
rect 491300 128 491352 134
rect 491300 70 491352 76
rect 492282 -960 492394 190
rect 492496 138 492548 144
rect 492588 196 492640 202
rect 492588 138 492640 144
rect 493478 -960 493590 326
rect 494674 -960 494786 480
rect 495544 354 495572 682
rect 495870 354 495982 480
rect 495544 326 495982 354
rect 495870 -960 495982 326
rect 496740 66 496768 3060
rect 497096 808 497148 814
rect 497096 750 497148 756
rect 497108 480 497136 750
rect 496728 60 496780 66
rect 496728 2 496780 8
rect 497066 -960 497178 480
rect 497936 406 497964 3060
rect 498936 876 498988 882
rect 498936 818 498988 824
rect 498200 604 498252 610
rect 498200 546 498252 552
rect 498212 480 498240 546
rect 497924 400 497976 406
rect 497924 342 497976 348
rect 498170 -960 498282 480
rect 498948 354 498976 818
rect 499040 814 499068 3060
rect 499028 808 499080 814
rect 499028 750 499080 756
rect 499366 354 499478 480
rect 500144 474 500172 3060
rect 501248 1222 501276 3060
rect 501236 1216 501288 1222
rect 501236 1158 501288 1164
rect 501420 1148 501472 1154
rect 501420 1090 501472 1096
rect 500592 672 500644 678
rect 500592 614 500644 620
rect 500604 480 500632 614
rect 500132 468 500184 474
rect 500132 410 500184 416
rect 498948 326 499478 354
rect 499366 -960 499478 326
rect 500562 -960 500674 480
rect 501432 354 501460 1090
rect 502260 746 502288 3060
rect 502984 1012 503036 1018
rect 502984 954 503036 960
rect 502248 740 502300 746
rect 502248 682 502300 688
rect 502996 480 503024 954
rect 503456 678 503484 3060
rect 503444 672 503496 678
rect 503444 614 503496 620
rect 503812 604 503864 610
rect 503812 546 503864 552
rect 501758 354 501870 480
rect 501432 326 501870 354
rect 501758 -960 501870 326
rect 502954 -960 503066 480
rect 503824 354 503852 546
rect 504150 354 504262 480
rect 504560 406 504588 3060
rect 503824 326 504262 354
rect 504548 400 504600 406
rect 504548 342 504600 348
rect 504150 -960 504262 326
rect 505346 82 505458 480
rect 505664 338 505692 3060
rect 506768 1154 506796 3060
rect 507780 1290 507808 3060
rect 507308 1284 507360 1290
rect 507308 1226 507360 1232
rect 507768 1284 507820 1290
rect 507768 1226 507820 1232
rect 506756 1148 506808 1154
rect 506756 1090 506808 1096
rect 505652 332 505704 338
rect 505652 274 505704 280
rect 506450 218 506562 480
rect 507320 354 507348 1226
rect 508872 944 508924 950
rect 508872 886 508924 892
rect 508884 480 508912 886
rect 508976 610 509004 3060
rect 510080 1358 510108 3060
rect 511198 3046 511488 3074
rect 512302 3046 512684 3074
rect 509700 1352 509752 1358
rect 509700 1294 509752 1300
rect 510068 1352 510120 1358
rect 510068 1294 510120 1300
rect 508964 604 509016 610
rect 508964 546 509016 552
rect 507646 354 507758 480
rect 507320 326 507758 354
rect 506450 202 506704 218
rect 506450 196 506716 202
rect 506450 190 506664 196
rect 505560 128 505612 134
rect 505346 76 505560 82
rect 505346 70 505612 76
rect 505346 54 505600 70
rect 505346 -960 505458 54
rect 506450 -960 506562 190
rect 506664 138 506716 144
rect 507646 -960 507758 326
rect 508842 -960 508954 480
rect 509712 354 509740 1294
rect 510038 354 510150 480
rect 509712 326 510150 354
rect 510038 -960 510150 326
rect 511234 82 511346 480
rect 511460 270 511488 3046
rect 512092 536 512144 542
rect 512092 478 512144 484
rect 512104 354 512132 478
rect 512430 354 512542 480
rect 512104 326 512542 354
rect 511448 264 511500 270
rect 511448 206 511500 212
rect 511234 66 511488 82
rect 511234 60 511500 66
rect 511234 54 511448 60
rect 511234 -960 511346 54
rect 511448 2 511500 8
rect 512430 -960 512542 326
rect 512656 202 512684 3046
rect 513300 2990 513328 3060
rect 513288 2984 513340 2990
rect 513288 2926 513340 2932
rect 513564 808 513616 814
rect 513564 750 513616 756
rect 513576 480 513604 750
rect 512644 196 512696 202
rect 512644 138 512696 144
rect 513534 -960 513646 480
rect 514496 134 514524 3060
rect 515496 1216 515548 1222
rect 515496 1158 515548 1164
rect 514730 354 514842 480
rect 514944 468 514996 474
rect 514944 410 514996 416
rect 514956 354 514984 410
rect 514730 326 514984 354
rect 515508 354 515536 1158
rect 515600 950 515628 3060
rect 516704 1222 516732 3060
rect 517520 2916 517572 2922
rect 517520 2858 517572 2864
rect 517532 1290 517560 2858
rect 517612 2848 517664 2854
rect 517612 2790 517664 2796
rect 517520 1284 517572 1290
rect 517520 1226 517572 1232
rect 516692 1216 516744 1222
rect 516692 1158 516744 1164
rect 517624 1154 517652 2790
rect 517612 1148 517664 1154
rect 517612 1090 517664 1096
rect 515588 944 515640 950
rect 515588 886 515640 892
rect 517152 740 517204 746
rect 517152 682 517204 688
rect 517164 480 517192 682
rect 517808 542 517836 3060
rect 518820 1086 518848 3060
rect 518808 1080 518860 1086
rect 518808 1022 518860 1028
rect 520016 1018 520044 3060
rect 520004 1012 520056 1018
rect 520004 954 520056 960
rect 521120 746 521148 3060
rect 521844 2848 521896 2854
rect 521844 2790 521896 2796
rect 521108 740 521160 746
rect 521108 682 521160 688
rect 518348 672 518400 678
rect 518348 614 518400 620
rect 517796 536 517848 542
rect 515926 354 516038 480
rect 515508 326 516038 354
rect 514484 128 514536 134
rect 514484 70 514536 76
rect 514730 -960 514842 326
rect 515926 -960 516038 326
rect 517122 -960 517234 480
rect 517796 478 517848 484
rect 518360 480 518388 614
rect 521856 480 521884 2790
rect 522224 1154 522252 3060
rect 523040 2916 523092 2922
rect 523040 2858 523092 2864
rect 522212 1148 522264 1154
rect 522212 1090 522264 1096
rect 523052 480 523080 2858
rect 523328 678 523356 3060
rect 524340 678 524368 3060
rect 525550 3046 525748 3074
rect 526654 3046 526944 3074
rect 525432 1352 525484 1358
rect 525432 1294 525484 1300
rect 523316 672 523368 678
rect 523316 614 523368 620
rect 524328 672 524380 678
rect 524328 614 524380 620
rect 523868 604 523920 610
rect 523868 546 523920 552
rect 518318 -960 518430 480
rect 519514 354 519626 480
rect 519728 400 519780 406
rect 519514 348 519728 354
rect 520710 354 520822 480
rect 519514 342 519780 348
rect 519514 326 519768 342
rect 520384 338 520822 354
rect 520372 332 520822 338
rect 519514 -960 519626 326
rect 520424 326 520822 332
rect 520372 274 520424 280
rect 520710 -960 520822 326
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 523880 354 523908 546
rect 525444 480 525472 1294
rect 524206 354 524318 480
rect 523880 326 524318 354
rect 524206 -960 524318 326
rect 525402 -960 525514 480
rect 525720 474 525748 3046
rect 525800 2916 525852 2922
rect 525800 2858 525852 2864
rect 525812 950 525840 2858
rect 525800 944 525852 950
rect 525800 886 525852 892
rect 525708 468 525760 474
rect 525708 410 525760 416
rect 526260 264 526312 270
rect 526598 218 526710 480
rect 526312 212 526710 218
rect 526260 206 526710 212
rect 526272 190 526710 206
rect 526598 -960 526710 190
rect 526916 66 526944 3046
rect 527744 882 527772 3060
rect 527732 876 527784 882
rect 527732 818 527784 824
rect 528848 814 528876 3060
rect 529966 3058 530072 3074
rect 529966 3052 530084 3058
rect 529966 3046 530032 3052
rect 530032 2994 530084 3000
rect 529020 2984 529072 2990
rect 529020 2926 529072 2932
rect 528836 808 528888 814
rect 528836 750 528888 756
rect 529032 480 529060 2926
rect 527794 218 527906 480
rect 527794 202 528048 218
rect 527794 196 528060 202
rect 527794 190 528008 196
rect 526904 60 526956 66
rect 526904 2 526956 8
rect 527794 -960 527906 190
rect 528008 138 528060 144
rect 528990 -960 529102 480
rect 529940 128 529992 134
rect 530094 82 530206 480
rect 531056 338 531084 3060
rect 531320 2916 531372 2922
rect 531320 2858 531372 2864
rect 531332 480 531360 2858
rect 532056 1216 532108 1222
rect 532056 1158 532108 1164
rect 531044 332 531096 338
rect 531044 274 531096 280
rect 529992 76 530206 82
rect 529940 70 530206 76
rect 529952 54 530206 70
rect 530094 -960 530206 54
rect 531290 -960 531402 480
rect 532068 354 532096 1158
rect 532160 950 532188 3060
rect 533278 3046 533844 3074
rect 543214 3068 543464 3074
rect 560484 3120 560536 3126
rect 543214 3062 543516 3068
rect 532148 944 532200 950
rect 532148 886 532200 892
rect 533252 672 533304 678
rect 533252 614 533304 620
rect 532486 354 532598 480
rect 533264 406 533292 614
rect 533816 610 533844 3046
rect 534368 1290 534396 3060
rect 534356 1284 534408 1290
rect 534356 1226 534408 1232
rect 534540 1080 534592 1086
rect 534540 1022 534592 1028
rect 533712 604 533764 610
rect 533712 546 533764 552
rect 533804 604 533856 610
rect 533804 546 533856 552
rect 533724 480 533752 546
rect 532068 326 532598 354
rect 533252 400 533304 406
rect 533252 342 533304 348
rect 532486 -960 532598 326
rect 533682 -960 533794 480
rect 534552 354 534580 1022
rect 534878 354 534990 480
rect 534552 326 534990 354
rect 534878 -960 534990 326
rect 535380 202 535408 3060
rect 536576 2922 536604 3060
rect 536564 2916 536616 2922
rect 536564 2858 536616 2864
rect 536104 1012 536156 1018
rect 536104 954 536156 960
rect 536116 480 536144 954
rect 537680 746 537708 3060
rect 538128 1148 538180 1154
rect 538128 1090 538180 1096
rect 537208 740 537260 746
rect 537208 682 537260 688
rect 537668 740 537720 746
rect 537668 682 537720 688
rect 537220 480 537248 682
rect 535368 196 535420 202
rect 535368 138 535420 144
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538140 354 538168 1090
rect 538374 354 538486 480
rect 538140 326 538486 354
rect 538374 -960 538486 326
rect 538784 270 538812 3060
rect 539888 1358 539916 3060
rect 539876 1352 539928 1358
rect 539876 1294 539928 1300
rect 539600 672 539652 678
rect 539600 614 539652 620
rect 540900 626 540928 3060
rect 542096 678 542124 3060
rect 543214 3046 543504 3062
rect 544318 3046 544608 3074
rect 544384 876 544436 882
rect 544384 818 544436 824
rect 542084 672 542136 678
rect 539612 480 539640 614
rect 540900 598 541020 626
rect 542084 614 542136 620
rect 538772 264 538824 270
rect 538772 206 538824 212
rect 539570 -960 539682 480
rect 540428 400 540480 406
rect 540766 354 540878 480
rect 540480 348 540878 354
rect 540428 342 540878 348
rect 540440 326 540878 342
rect 540766 -960 540878 326
rect 540992 134 541020 598
rect 544396 480 544424 818
rect 541962 354 542074 480
rect 542176 468 542228 474
rect 542176 410 542228 416
rect 542188 354 542216 410
rect 541962 326 542216 354
rect 540980 128 541032 134
rect 540980 70 541032 76
rect 541962 -960 542074 326
rect 543158 82 543270 480
rect 542832 66 543270 82
rect 542820 60 543270 66
rect 542872 54 543270 60
rect 542820 2 542872 8
rect 543158 -960 543270 54
rect 544354 -960 544466 480
rect 544580 474 544608 3046
rect 545408 610 545436 3060
rect 545488 808 545540 814
rect 545488 750 545540 756
rect 545396 604 545448 610
rect 545396 546 545448 552
rect 545500 480 545528 750
rect 544568 468 544620 474
rect 544568 410 544620 416
rect 545458 -960 545570 480
rect 546420 66 546448 3060
rect 546684 3052 546736 3058
rect 546684 2994 546736 3000
rect 546696 480 546724 2994
rect 547616 882 547644 3060
rect 548734 3046 549024 3074
rect 548708 944 548760 950
rect 548708 886 548760 892
rect 547604 876 547656 882
rect 547604 818 547656 824
rect 546408 60 546460 66
rect 546408 2 546460 8
rect 546654 -960 546766 480
rect 547850 354 547962 480
rect 548720 354 548748 886
rect 548996 678 549024 3046
rect 549824 2990 549852 3060
rect 549812 2984 549864 2990
rect 549812 2926 549864 2932
rect 550928 814 550956 3060
rect 551100 1284 551152 1290
rect 551100 1226 551152 1232
rect 550916 808 550968 814
rect 550916 750 550968 756
rect 548984 672 549036 678
rect 548984 614 549036 620
rect 549046 354 549158 480
rect 547850 338 548104 354
rect 547850 332 548116 338
rect 547850 326 548064 332
rect 547850 -960 547962 326
rect 548720 326 549158 354
rect 548064 274 548116 280
rect 549046 -960 549158 326
rect 550242 354 550354 480
rect 550456 400 550508 406
rect 550242 348 550456 354
rect 550242 342 550508 348
rect 551112 354 551140 1226
rect 551438 354 551550 480
rect 550242 326 550496 342
rect 551112 326 551550 354
rect 551940 338 551968 3060
rect 553150 3058 553348 3074
rect 553150 3052 553360 3058
rect 553150 3046 553308 3052
rect 553308 2994 553360 3000
rect 553768 2916 553820 2922
rect 553768 2858 553820 2864
rect 553780 480 553808 2858
rect 550242 -960 550354 326
rect 551438 -960 551550 326
rect 551928 332 551980 338
rect 551928 274 551980 280
rect 552634 218 552746 480
rect 552634 202 552888 218
rect 552634 196 552900 202
rect 552634 190 552848 196
rect 552634 -960 552746 190
rect 552848 138 552900 144
rect 553738 -960 553850 480
rect 554240 202 554268 3060
rect 554964 740 555016 746
rect 554964 682 555016 688
rect 554976 480 555004 682
rect 554228 196 554280 202
rect 554228 138 554280 144
rect 554934 -960 555046 480
rect 555344 406 555372 3060
rect 557184 3046 557474 3074
rect 558670 3046 558868 3074
rect 562232 3120 562284 3126
rect 560484 3062 560536 3068
rect 561982 3068 562232 3074
rect 561982 3062 562284 3068
rect 556988 1352 557040 1358
rect 556988 1294 557040 1300
rect 555332 400 555384 406
rect 555332 342 555384 348
rect 556130 218 556242 480
rect 556344 264 556396 270
rect 556130 212 556344 218
rect 556130 206 556396 212
rect 556130 190 556384 206
rect 556130 -960 556242 190
rect 557000 82 557028 1294
rect 557184 270 557212 3046
rect 557172 264 557224 270
rect 557172 206 557224 212
rect 557326 82 557438 480
rect 557000 54 557438 82
rect 557326 -960 557438 54
rect 558522 82 558634 480
rect 558840 134 558868 3046
rect 559760 2922 559788 3060
rect 559748 2916 559800 2922
rect 559748 2858 559800 2864
rect 559380 536 559432 542
rect 559380 478 559432 484
rect 559392 354 559420 478
rect 559718 354 559830 480
rect 559392 326 559830 354
rect 560496 354 560524 3062
rect 561982 3046 562272 3062
rect 562980 2854 563008 3060
rect 571524 3052 571576 3058
rect 571524 2994 571576 3000
rect 568028 2984 568080 2990
rect 568028 2926 568080 2932
rect 562968 2848 563020 2854
rect 562968 2790 563020 2796
rect 565636 876 565688 882
rect 565636 818 565688 824
rect 563244 604 563296 610
rect 563244 546 563296 552
rect 563256 480 563284 546
rect 565648 480 565676 818
rect 566832 672 566884 678
rect 566832 614 566884 620
rect 566844 480 566872 614
rect 568040 480 568068 2926
rect 569132 808 569184 814
rect 569132 750 569184 756
rect 569144 480 569172 750
rect 571536 480 571564 2994
rect 575124 480 575152 3198
rect 579804 3188 579856 3194
rect 579804 3130 579856 3136
rect 578608 2916 578660 2922
rect 578608 2858 578660 2864
rect 578620 480 578648 2858
rect 579816 480 579844 3130
rect 581000 3120 581052 3126
rect 581000 3062 581052 3068
rect 581012 480 581040 3062
rect 582196 2848 582248 2854
rect 582196 2790 582248 2796
rect 582208 480 582236 2790
rect 583404 480 583432 3266
rect 560822 354 560934 480
rect 560496 326 560934 354
rect 558736 128 558788 134
rect 558522 76 558736 82
rect 558522 70 558788 76
rect 558828 128 558880 134
rect 558828 70 558880 76
rect 558522 54 558776 70
rect 558522 -960 558634 54
rect 559718 -960 559830 326
rect 560822 -960 560934 326
rect 562018 354 562130 480
rect 562232 468 562284 474
rect 562232 410 562284 416
rect 562244 354 562272 410
rect 562018 326 562272 354
rect 562018 -960 562130 326
rect 563214 -960 563326 480
rect 564410 82 564522 480
rect 564410 66 564664 82
rect 564410 60 564676 66
rect 564410 54 564624 60
rect 564410 -960 564522 54
rect 564624 2 564676 8
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 354 570410 480
rect 570298 338 570552 354
rect 570298 332 570564 338
rect 570298 326 570512 332
rect 570298 -960 570410 326
rect 570512 274 570564 280
rect 571494 -960 571606 480
rect 572690 218 572802 480
rect 573548 400 573600 406
rect 573886 354 573998 480
rect 573600 348 573998 354
rect 573548 342 573998 348
rect 573560 326 573998 342
rect 572690 202 572944 218
rect 572690 196 572956 202
rect 572690 190 572904 196
rect 572690 -960 572802 190
rect 572904 138 572956 144
rect 573886 -960 573998 326
rect 575082 -960 575194 480
rect 575940 264 575992 270
rect 576278 218 576390 480
rect 575992 212 576390 218
rect 575940 206 576390 212
rect 575952 190 576390 206
rect 576278 -960 576390 190
rect 577136 128 577188 134
rect 577382 82 577494 480
rect 577188 76 577494 82
rect 577136 70 577494 76
rect 577148 54 577494 70
rect 577382 -960 577494 54
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 2778 697312 2834 697368
rect 581642 697176 581698 697232
rect 581642 691464 581698 691520
rect 2778 690784 2834 690840
rect 2778 684256 2834 684312
rect 582378 683848 582434 683904
rect 582378 678408 582434 678464
rect 2778 678000 2834 678056
rect 2778 671200 2834 671256
rect 582378 670656 582434 670712
rect 582378 665352 582434 665408
rect 2778 665216 2834 665272
rect 2778 658144 2834 658200
rect 582378 657328 582434 657384
rect 2778 652432 2834 652488
rect 582378 652296 582434 652352
rect 2778 645088 2834 645144
rect 581642 644000 581698 644056
rect 2778 639648 2834 639704
rect 581642 639240 581698 639296
rect 2778 632032 2834 632088
rect 582378 630808 582434 630864
rect 2778 626864 2834 626920
rect 582378 626184 582434 626240
rect 2778 619112 2834 619168
rect 581642 617480 581698 617536
rect 2778 613944 2834 614000
rect 581642 613128 581698 613184
rect 2778 606056 2834 606112
rect 581642 604152 581698 604208
rect 2778 601296 2834 601352
rect 581642 600072 581698 600128
rect 1582 593000 1638 593056
rect 581642 590960 581698 591016
rect 1582 588512 1638 588568
rect 581642 587016 581698 587072
rect 2042 579944 2098 580000
rect 581642 577632 581698 577688
rect 2042 575728 2098 575784
rect 581642 573960 581698 574016
rect 1490 566888 1546 566944
rect 582378 564304 582434 564360
rect 1490 562944 1546 563000
rect 582378 560904 582434 560960
rect 1490 553832 1546 553888
rect 581642 551112 581698 551168
rect 1490 550160 1546 550216
rect 581642 547712 581698 547768
rect 1398 540776 1454 540832
rect 582378 537784 582434 537840
rect 1398 537376 1454 537432
rect 582378 534792 582434 534848
rect 1490 527856 1546 527912
rect 1490 524592 1546 524648
rect 582378 524456 582434 524512
rect 582378 521736 582434 521792
rect 1582 514800 1638 514856
rect 1582 511808 1638 511864
rect 582378 511264 582434 511320
rect 582378 508680 582434 508736
rect 1582 501744 1638 501800
rect 1582 499024 1638 499080
rect 581642 497936 581698 497992
rect 581642 495624 581698 495680
rect 1582 488688 1638 488744
rect 1582 486240 1638 486296
rect 582378 484608 582434 484664
rect 582378 482568 582434 482624
rect 2778 475632 2834 475688
rect 2778 473456 2834 473512
rect 581642 471416 581698 471472
rect 581642 469512 581698 469568
rect 1582 462576 1638 462632
rect 1582 460672 1638 460728
rect 581642 458088 581698 458144
rect 581642 456456 581698 456512
rect 2778 449520 2834 449576
rect 2778 447888 2834 447944
rect 2778 436600 2834 436656
rect 2778 435104 2834 435160
rect 2778 423544 2834 423600
rect 2778 422320 2834 422376
rect 1306 294344 1362 294400
rect 1306 293120 1362 293176
rect 2778 281560 2834 281616
rect 2778 280064 2834 280120
rect 1306 268776 1362 268832
rect 1306 267144 1362 267200
rect 582378 260480 582434 260536
rect 582378 258848 582434 258904
rect 1306 255992 1362 256048
rect 1306 254088 1362 254144
rect 580906 247016 580962 247072
rect 580906 245520 580962 245576
rect 2778 243208 2834 243264
rect 2778 241032 2834 241088
rect 582378 234368 582434 234424
rect 582378 232328 582434 232384
rect 2778 230560 2834 230616
rect 2778 227976 2834 228032
rect 580906 220904 580962 220960
rect 580906 219000 580962 219056
rect 2778 217640 2834 217696
rect 2778 214920 2834 214976
rect 582378 208256 582434 208312
rect 582378 205672 582434 205728
rect 2778 204856 2834 204912
rect 2778 201864 2834 201920
rect 580906 194656 580962 194712
rect 580906 192480 580962 192536
rect 1306 192072 1362 192128
rect 1306 188808 1362 188864
rect 580906 182416 580962 182472
rect 2778 179288 2834 179344
rect 580906 179152 580962 179208
rect 2778 175888 2834 175944
rect 580906 168544 580962 168600
rect 2778 166504 2834 166560
rect 580906 165824 580962 165880
rect 2778 162832 2834 162888
rect 580906 156304 580962 156360
rect 1306 153720 1362 153776
rect 580906 152632 580962 152688
rect 1306 149776 1362 149832
rect 580906 142568 580962 142624
rect 570 140936 626 140992
rect 580906 139304 580962 139360
rect 570 136720 626 136776
rect 580906 130192 580962 130248
rect 754 128152 810 128208
rect 580906 125976 580962 126032
rect 754 123664 810 123720
rect 579894 116320 579950 116376
rect 1306 115368 1362 115424
rect 579894 112784 579950 112840
rect 1306 110608 1362 110664
rect 580906 103536 580962 103592
rect 1582 102584 1638 102640
rect 580906 99456 580962 99512
rect 1582 97552 1638 97608
rect 580906 90208 580962 90264
rect 1582 89800 1638 89856
rect 580906 86128 580962 86184
rect 1582 84632 1638 84688
rect 579894 77288 579950 77344
rect 1582 77016 1638 77072
rect 579894 72936 579950 72992
rect 1582 71576 1638 71632
rect 1490 64232 1546 64288
rect 580906 64096 580962 64152
rect 580906 59608 580962 59664
rect 1490 58520 1546 58576
rect 2042 51448 2098 51504
rect 580906 51040 580962 51096
rect 580906 46280 580962 46336
rect 2042 45464 2098 45520
rect 2042 38664 2098 38720
rect 580906 37984 580962 38040
rect 580906 33088 580962 33144
rect 2042 32408 2098 32464
rect 1490 25880 1546 25936
rect 580906 24928 580962 24984
rect 580906 19760 580962 19816
rect 1490 19352 1546 19408
rect 2042 13096 2098 13152
rect 579894 12688 579950 12744
rect 579894 6568 579950 6624
rect 2042 6432 2098 6488
rect 70214 3884 70216 3904
rect 70216 3884 70268 3904
rect 70268 3884 70270 3904
rect 70214 3848 70270 3884
rect 73618 3848 73674 3904
rect 5446 312 5502 368
rect 6274 40 6330 96
rect 12162 448 12218 504
rect 13726 176 13782 232
rect 23938 312 23994 368
rect 25042 40 25098 96
rect 25686 312 25742 368
rect 28906 584 28962 640
rect 30838 448 30894 504
rect 31942 176 31998 232
rect 37002 176 37058 232
rect 42706 312 42762 368
rect 46294 584 46350 640
rect 46846 40 46902 96
rect 54022 176 54078 232
rect 62854 40 62910 96
<< metal3 >>
rect -960 697370 480 697460
rect 2773 697370 2839 697373
rect -960 697368 2839 697370
rect -960 697312 2778 697368
rect 2834 697312 2839 697368
rect -960 697310 2839 697312
rect -960 697220 480 697310
rect 2773 697307 2839 697310
rect 581637 697234 581703 697237
rect 583520 697234 584960 697324
rect 581637 697232 584960 697234
rect 581637 697176 581642 697232
rect 581698 697176 584960 697232
rect 581637 697174 584960 697176
rect 581637 697171 581703 697174
rect 583520 697084 584960 697174
rect 581637 691522 581703 691525
rect 580796 691520 581703 691522
rect 580796 691464 581642 691520
rect 581698 691464 581703 691520
rect 580796 691462 581703 691464
rect 581637 691459 581703 691462
rect 2773 690842 2839 690845
rect 2773 690840 3220 690842
rect 2773 690784 2778 690840
rect 2834 690784 3220 690840
rect 2773 690782 3220 690784
rect 2773 690779 2839 690782
rect -960 684314 480 684404
rect 2773 684314 2839 684317
rect -960 684312 2839 684314
rect -960 684256 2778 684312
rect 2834 684256 2839 684312
rect -960 684254 2839 684256
rect -960 684164 480 684254
rect 2773 684251 2839 684254
rect 582373 683906 582439 683909
rect 583520 683906 584960 683996
rect 582373 683904 584960 683906
rect 582373 683848 582378 683904
rect 582434 683848 584960 683904
rect 582373 683846 584960 683848
rect 582373 683843 582439 683846
rect 583520 683756 584960 683846
rect 582373 678466 582439 678469
rect 580796 678464 582439 678466
rect 580796 678408 582378 678464
rect 582434 678408 582439 678464
rect 580796 678406 582439 678408
rect 582373 678403 582439 678406
rect 2773 678058 2839 678061
rect 2773 678056 3220 678058
rect 2773 678000 2778 678056
rect 2834 678000 3220 678056
rect 2773 677998 3220 678000
rect 2773 677995 2839 677998
rect -960 671258 480 671348
rect 2773 671258 2839 671261
rect -960 671256 2839 671258
rect -960 671200 2778 671256
rect 2834 671200 2839 671256
rect -960 671198 2839 671200
rect -960 671108 480 671198
rect 2773 671195 2839 671198
rect 582373 670714 582439 670717
rect 583520 670714 584960 670804
rect 582373 670712 584960 670714
rect 582373 670656 582378 670712
rect 582434 670656 584960 670712
rect 582373 670654 584960 670656
rect 582373 670651 582439 670654
rect 583520 670564 584960 670654
rect 582373 665410 582439 665413
rect 580796 665408 582439 665410
rect 580796 665352 582378 665408
rect 582434 665352 582439 665408
rect 580796 665350 582439 665352
rect 582373 665347 582439 665350
rect 2773 665274 2839 665277
rect 2773 665272 3220 665274
rect 2773 665216 2778 665272
rect 2834 665216 3220 665272
rect 2773 665214 3220 665216
rect 2773 665211 2839 665214
rect -960 658202 480 658292
rect 2773 658202 2839 658205
rect -960 658200 2839 658202
rect -960 658144 2778 658200
rect 2834 658144 2839 658200
rect -960 658142 2839 658144
rect -960 658052 480 658142
rect 2773 658139 2839 658142
rect 582373 657386 582439 657389
rect 583520 657386 584960 657476
rect 582373 657384 584960 657386
rect 582373 657328 582378 657384
rect 582434 657328 584960 657384
rect 582373 657326 584960 657328
rect 582373 657323 582439 657326
rect 583520 657236 584960 657326
rect 2773 652490 2839 652493
rect 2773 652488 3220 652490
rect 2773 652432 2778 652488
rect 2834 652432 3220 652488
rect 2773 652430 3220 652432
rect 2773 652427 2839 652430
rect 582373 652354 582439 652357
rect 580796 652352 582439 652354
rect 580796 652296 582378 652352
rect 582434 652296 582439 652352
rect 580796 652294 582439 652296
rect 582373 652291 582439 652294
rect -960 645146 480 645236
rect 2773 645146 2839 645149
rect -960 645144 2839 645146
rect -960 645088 2778 645144
rect 2834 645088 2839 645144
rect -960 645086 2839 645088
rect -960 644996 480 645086
rect 2773 645083 2839 645086
rect 581637 644058 581703 644061
rect 583520 644058 584960 644148
rect 581637 644056 584960 644058
rect 581637 644000 581642 644056
rect 581698 644000 584960 644056
rect 581637 643998 584960 644000
rect 581637 643995 581703 643998
rect 583520 643908 584960 643998
rect 2773 639706 2839 639709
rect 2773 639704 3220 639706
rect 2773 639648 2778 639704
rect 2834 639648 3220 639704
rect 2773 639646 3220 639648
rect 2773 639643 2839 639646
rect 581637 639298 581703 639301
rect 580796 639296 581703 639298
rect 580796 639240 581642 639296
rect 581698 639240 581703 639296
rect 580796 639238 581703 639240
rect 581637 639235 581703 639238
rect -960 632090 480 632180
rect 2773 632090 2839 632093
rect -960 632088 2839 632090
rect -960 632032 2778 632088
rect 2834 632032 2839 632088
rect -960 632030 2839 632032
rect -960 631940 480 632030
rect 2773 632027 2839 632030
rect 582373 630866 582439 630869
rect 583520 630866 584960 630956
rect 582373 630864 584960 630866
rect 582373 630808 582378 630864
rect 582434 630808 584960 630864
rect 582373 630806 584960 630808
rect 582373 630803 582439 630806
rect 583520 630716 584960 630806
rect 2773 626922 2839 626925
rect 2773 626920 3220 626922
rect 2773 626864 2778 626920
rect 2834 626864 3220 626920
rect 2773 626862 3220 626864
rect 2773 626859 2839 626862
rect 582373 626242 582439 626245
rect 580796 626240 582439 626242
rect 580796 626184 582378 626240
rect 582434 626184 582439 626240
rect 580796 626182 582439 626184
rect 582373 626179 582439 626182
rect -960 619170 480 619260
rect 2773 619170 2839 619173
rect -960 619168 2839 619170
rect -960 619112 2778 619168
rect 2834 619112 2839 619168
rect -960 619110 2839 619112
rect -960 619020 480 619110
rect 2773 619107 2839 619110
rect 581637 617538 581703 617541
rect 583520 617538 584960 617628
rect 581637 617536 584960 617538
rect 581637 617480 581642 617536
rect 581698 617480 584960 617536
rect 581637 617478 584960 617480
rect 581637 617475 581703 617478
rect 583520 617388 584960 617478
rect 2773 614002 2839 614005
rect 2773 614000 3220 614002
rect 2773 613944 2778 614000
rect 2834 613944 3220 614000
rect 2773 613942 3220 613944
rect 2773 613939 2839 613942
rect 581637 613186 581703 613189
rect 580796 613184 581703 613186
rect 580796 613128 581642 613184
rect 581698 613128 581703 613184
rect 580796 613126 581703 613128
rect 581637 613123 581703 613126
rect -960 606114 480 606204
rect 2773 606114 2839 606117
rect -960 606112 2839 606114
rect -960 606056 2778 606112
rect 2834 606056 2839 606112
rect -960 606054 2839 606056
rect -960 605964 480 606054
rect 2773 606051 2839 606054
rect 581637 604210 581703 604213
rect 583520 604210 584960 604300
rect 581637 604208 584960 604210
rect 581637 604152 581642 604208
rect 581698 604152 584960 604208
rect 581637 604150 584960 604152
rect 581637 604147 581703 604150
rect 583520 604060 584960 604150
rect 2773 601354 2839 601357
rect 2773 601352 3220 601354
rect 2773 601296 2778 601352
rect 2834 601296 3220 601352
rect 2773 601294 3220 601296
rect 2773 601291 2839 601294
rect 581637 600130 581703 600133
rect 580796 600128 581703 600130
rect 580796 600072 581642 600128
rect 581698 600072 581703 600128
rect 580796 600070 581703 600072
rect 581637 600067 581703 600070
rect -960 593058 480 593148
rect 1577 593058 1643 593061
rect -960 593056 1643 593058
rect -960 593000 1582 593056
rect 1638 593000 1643 593056
rect -960 592998 1643 593000
rect -960 592908 480 592998
rect 1577 592995 1643 592998
rect 581637 591018 581703 591021
rect 583520 591018 584960 591108
rect 581637 591016 584960 591018
rect 581637 590960 581642 591016
rect 581698 590960 584960 591016
rect 581637 590958 584960 590960
rect 581637 590955 581703 590958
rect 583520 590868 584960 590958
rect 1577 588570 1643 588573
rect 1577 588568 3220 588570
rect 1577 588512 1582 588568
rect 1638 588512 3220 588568
rect 1577 588510 3220 588512
rect 1577 588507 1643 588510
rect 581637 587074 581703 587077
rect 580796 587072 581703 587074
rect 580796 587016 581642 587072
rect 581698 587016 581703 587072
rect 580796 587014 581703 587016
rect 581637 587011 581703 587014
rect -960 580002 480 580092
rect 2037 580002 2103 580005
rect -960 580000 2103 580002
rect -960 579944 2042 580000
rect 2098 579944 2103 580000
rect -960 579942 2103 579944
rect -960 579852 480 579942
rect 2037 579939 2103 579942
rect 581637 577690 581703 577693
rect 583520 577690 584960 577780
rect 581637 577688 584960 577690
rect 581637 577632 581642 577688
rect 581698 577632 584960 577688
rect 581637 577630 584960 577632
rect 581637 577627 581703 577630
rect 583520 577540 584960 577630
rect 2037 575786 2103 575789
rect 2037 575784 3220 575786
rect 2037 575728 2042 575784
rect 2098 575728 3220 575784
rect 2037 575726 3220 575728
rect 2037 575723 2103 575726
rect 581637 574018 581703 574021
rect 580796 574016 581703 574018
rect 580796 573960 581642 574016
rect 581698 573960 581703 574016
rect 580796 573958 581703 573960
rect 581637 573955 581703 573958
rect -960 566946 480 567036
rect 1485 566946 1551 566949
rect -960 566944 1551 566946
rect -960 566888 1490 566944
rect 1546 566888 1551 566944
rect -960 566886 1551 566888
rect -960 566796 480 566886
rect 1485 566883 1551 566886
rect 582373 564362 582439 564365
rect 583520 564362 584960 564452
rect 582373 564360 584960 564362
rect 582373 564304 582378 564360
rect 582434 564304 584960 564360
rect 582373 564302 584960 564304
rect 582373 564299 582439 564302
rect 583520 564212 584960 564302
rect 1485 563002 1551 563005
rect 1485 563000 3220 563002
rect 1485 562944 1490 563000
rect 1546 562944 3220 563000
rect 1485 562942 3220 562944
rect 1485 562939 1551 562942
rect 582373 560962 582439 560965
rect 580796 560960 582439 560962
rect 580796 560904 582378 560960
rect 582434 560904 582439 560960
rect 580796 560902 582439 560904
rect 582373 560899 582439 560902
rect -960 553890 480 553980
rect 1485 553890 1551 553893
rect -960 553888 1551 553890
rect -960 553832 1490 553888
rect 1546 553832 1551 553888
rect -960 553830 1551 553832
rect -960 553740 480 553830
rect 1485 553827 1551 553830
rect 581637 551170 581703 551173
rect 583520 551170 584960 551260
rect 581637 551168 584960 551170
rect 581637 551112 581642 551168
rect 581698 551112 584960 551168
rect 581637 551110 584960 551112
rect 581637 551107 581703 551110
rect 583520 551020 584960 551110
rect 1485 550218 1551 550221
rect 1485 550216 3220 550218
rect 1485 550160 1490 550216
rect 1546 550160 3220 550216
rect 1485 550158 3220 550160
rect 1485 550155 1551 550158
rect 581637 547770 581703 547773
rect 580796 547768 581703 547770
rect 580796 547712 581642 547768
rect 581698 547712 581703 547768
rect 580796 547710 581703 547712
rect 581637 547707 581703 547710
rect -960 540834 480 540924
rect 1393 540834 1459 540837
rect -960 540832 1459 540834
rect -960 540776 1398 540832
rect 1454 540776 1459 540832
rect -960 540774 1459 540776
rect -960 540684 480 540774
rect 1393 540771 1459 540774
rect 582373 537842 582439 537845
rect 583520 537842 584960 537932
rect 582373 537840 584960 537842
rect 582373 537784 582378 537840
rect 582434 537784 584960 537840
rect 582373 537782 584960 537784
rect 582373 537779 582439 537782
rect 583520 537692 584960 537782
rect 1393 537434 1459 537437
rect 1393 537432 3220 537434
rect 1393 537376 1398 537432
rect 1454 537376 3220 537432
rect 1393 537374 3220 537376
rect 1393 537371 1459 537374
rect 582373 534850 582439 534853
rect 580796 534848 582439 534850
rect 580796 534792 582378 534848
rect 582434 534792 582439 534848
rect 580796 534790 582439 534792
rect 582373 534787 582439 534790
rect -960 527914 480 528004
rect 1485 527914 1551 527917
rect -960 527912 1551 527914
rect -960 527856 1490 527912
rect 1546 527856 1551 527912
rect -960 527854 1551 527856
rect -960 527764 480 527854
rect 1485 527851 1551 527854
rect 1485 524650 1551 524653
rect 1485 524648 3220 524650
rect 1485 524592 1490 524648
rect 1546 524592 3220 524648
rect 1485 524590 3220 524592
rect 1485 524587 1551 524590
rect 582373 524514 582439 524517
rect 583520 524514 584960 524604
rect 582373 524512 584960 524514
rect 582373 524456 582378 524512
rect 582434 524456 584960 524512
rect 582373 524454 584960 524456
rect 582373 524451 582439 524454
rect 583520 524364 584960 524454
rect 582373 521794 582439 521797
rect 580796 521792 582439 521794
rect 580796 521736 582378 521792
rect 582434 521736 582439 521792
rect 580796 521734 582439 521736
rect 582373 521731 582439 521734
rect -960 514858 480 514948
rect 1577 514858 1643 514861
rect -960 514856 1643 514858
rect -960 514800 1582 514856
rect 1638 514800 1643 514856
rect -960 514798 1643 514800
rect -960 514708 480 514798
rect 1577 514795 1643 514798
rect 1577 511866 1643 511869
rect 1577 511864 3220 511866
rect 1577 511808 1582 511864
rect 1638 511808 3220 511864
rect 1577 511806 3220 511808
rect 1577 511803 1643 511806
rect 582373 511322 582439 511325
rect 583520 511322 584960 511412
rect 582373 511320 584960 511322
rect 582373 511264 582378 511320
rect 582434 511264 584960 511320
rect 582373 511262 584960 511264
rect 582373 511259 582439 511262
rect 583520 511172 584960 511262
rect 582373 508738 582439 508741
rect 580796 508736 582439 508738
rect 580796 508680 582378 508736
rect 582434 508680 582439 508736
rect 580796 508678 582439 508680
rect 582373 508675 582439 508678
rect -960 501802 480 501892
rect 1577 501802 1643 501805
rect -960 501800 1643 501802
rect -960 501744 1582 501800
rect 1638 501744 1643 501800
rect -960 501742 1643 501744
rect -960 501652 480 501742
rect 1577 501739 1643 501742
rect 1577 499082 1643 499085
rect 1577 499080 3220 499082
rect 1577 499024 1582 499080
rect 1638 499024 3220 499080
rect 1577 499022 3220 499024
rect 1577 499019 1643 499022
rect 581637 497994 581703 497997
rect 583520 497994 584960 498084
rect 581637 497992 584960 497994
rect 581637 497936 581642 497992
rect 581698 497936 584960 497992
rect 581637 497934 584960 497936
rect 581637 497931 581703 497934
rect 583520 497844 584960 497934
rect 581637 495682 581703 495685
rect 580796 495680 581703 495682
rect 580796 495624 581642 495680
rect 581698 495624 581703 495680
rect 580796 495622 581703 495624
rect 581637 495619 581703 495622
rect -960 488746 480 488836
rect 1577 488746 1643 488749
rect -960 488744 1643 488746
rect -960 488688 1582 488744
rect 1638 488688 1643 488744
rect -960 488686 1643 488688
rect -960 488596 480 488686
rect 1577 488683 1643 488686
rect 1577 486298 1643 486301
rect 1577 486296 3220 486298
rect 1577 486240 1582 486296
rect 1638 486240 3220 486296
rect 1577 486238 3220 486240
rect 1577 486235 1643 486238
rect 582373 484666 582439 484669
rect 583520 484666 584960 484756
rect 582373 484664 584960 484666
rect 582373 484608 582378 484664
rect 582434 484608 584960 484664
rect 582373 484606 584960 484608
rect 582373 484603 582439 484606
rect 583520 484516 584960 484606
rect 582373 482626 582439 482629
rect 580796 482624 582439 482626
rect 580796 482568 582378 482624
rect 582434 482568 582439 482624
rect 580796 482566 582439 482568
rect 582373 482563 582439 482566
rect -960 475690 480 475780
rect 2773 475690 2839 475693
rect -960 475688 2839 475690
rect -960 475632 2778 475688
rect 2834 475632 2839 475688
rect -960 475630 2839 475632
rect -960 475540 480 475630
rect 2773 475627 2839 475630
rect 2773 473514 2839 473517
rect 2773 473512 3220 473514
rect 2773 473456 2778 473512
rect 2834 473456 3220 473512
rect 2773 473454 3220 473456
rect 2773 473451 2839 473454
rect 581637 471474 581703 471477
rect 583520 471474 584960 471564
rect 581637 471472 584960 471474
rect 581637 471416 581642 471472
rect 581698 471416 584960 471472
rect 581637 471414 584960 471416
rect 581637 471411 581703 471414
rect 583520 471324 584960 471414
rect 581637 469570 581703 469573
rect 580796 469568 581703 469570
rect 580796 469512 581642 469568
rect 581698 469512 581703 469568
rect 580796 469510 581703 469512
rect 581637 469507 581703 469510
rect -960 462634 480 462724
rect 1577 462634 1643 462637
rect -960 462632 1643 462634
rect -960 462576 1582 462632
rect 1638 462576 1643 462632
rect -960 462574 1643 462576
rect -960 462484 480 462574
rect 1577 462571 1643 462574
rect 1577 460730 1643 460733
rect 1577 460728 3220 460730
rect 1577 460672 1582 460728
rect 1638 460672 3220 460728
rect 1577 460670 3220 460672
rect 1577 460667 1643 460670
rect 581637 458146 581703 458149
rect 583520 458146 584960 458236
rect 581637 458144 584960 458146
rect 581637 458088 581642 458144
rect 581698 458088 584960 458144
rect 581637 458086 584960 458088
rect 581637 458083 581703 458086
rect 583520 457996 584960 458086
rect 581637 456514 581703 456517
rect 580796 456512 581703 456514
rect 580796 456456 581642 456512
rect 581698 456456 581703 456512
rect 580796 456454 581703 456456
rect 581637 456451 581703 456454
rect -960 449578 480 449668
rect 2773 449578 2839 449581
rect -960 449576 2839 449578
rect -960 449520 2778 449576
rect 2834 449520 2839 449576
rect -960 449518 2839 449520
rect -960 449428 480 449518
rect 2773 449515 2839 449518
rect 2773 447946 2839 447949
rect 2773 447944 3220 447946
rect 2773 447888 2778 447944
rect 2834 447888 3220 447944
rect 2773 447886 3220 447888
rect 2773 447883 2839 447886
rect 583520 444818 584960 444908
rect 583342 444758 584960 444818
rect 583342 444682 583402 444758
rect 583520 444682 584960 444758
rect 583342 444668 584960 444682
rect 583342 444622 583586 444668
rect 583526 444138 583586 444622
rect 580766 444078 583586 444138
rect 580766 443428 580826 444078
rect -960 436658 480 436748
rect 2773 436658 2839 436661
rect -960 436656 2839 436658
rect -960 436600 2778 436656
rect 2834 436600 2839 436656
rect -960 436598 2839 436600
rect -960 436508 480 436598
rect 2773 436595 2839 436598
rect 2773 435162 2839 435165
rect 2773 435160 3220 435162
rect 2773 435104 2778 435160
rect 2834 435104 3220 435160
rect 2773 435102 3220 435104
rect 2773 435099 2839 435102
rect 583520 431626 584960 431716
rect 583342 431566 584960 431626
rect 583342 431490 583402 431566
rect 583520 431490 584960 431566
rect 583342 431476 584960 431490
rect 583342 431430 583586 431476
rect 583526 431082 583586 431430
rect 580766 431022 583586 431082
rect 580766 430372 580826 431022
rect -960 423602 480 423692
rect 2773 423602 2839 423605
rect -960 423600 2839 423602
rect -960 423544 2778 423600
rect 2834 423544 2839 423600
rect -960 423542 2839 423544
rect -960 423452 480 423542
rect 2773 423539 2839 423542
rect 2773 422378 2839 422381
rect 2773 422376 3220 422378
rect 2773 422320 2778 422376
rect 2834 422320 3220 422376
rect 2773 422318 3220 422320
rect 2773 422315 2839 422318
rect 583520 418298 584960 418388
rect 583342 418238 584960 418298
rect 583342 418162 583402 418238
rect 583520 418162 584960 418238
rect 583342 418148 584960 418162
rect 583342 418102 583586 418148
rect 583526 417754 583586 418102
rect 580766 417694 583586 417754
rect 580766 417316 580826 417694
rect -960 410546 480 410636
rect -960 410486 3250 410546
rect -960 410396 480 410486
rect 3190 409564 3250 410486
rect 583520 404970 584960 405060
rect 580766 404910 584960 404970
rect 580766 404260 580826 404910
rect 583520 404820 584960 404910
rect -960 397490 480 397580
rect -960 397430 3250 397490
rect -960 397340 480 397430
rect 3190 396780 3250 397430
rect 583520 391778 584960 391868
rect 580766 391718 584960 391778
rect 580766 391204 580826 391718
rect 583520 391628 584960 391718
rect -960 384434 480 384524
rect -960 384374 3250 384434
rect -960 384284 480 384374
rect 3190 383996 3250 384374
rect 583520 378450 584960 378540
rect 580766 378390 584960 378450
rect 580766 378148 580826 378390
rect 583520 378300 584960 378390
rect -960 371378 480 371468
rect -960 371318 3250 371378
rect -960 371228 480 371318
rect 3190 371212 3250 371318
rect 583520 365122 584960 365212
rect 580796 365062 584960 365122
rect 583520 364972 584960 365062
rect -960 358458 480 358548
rect -960 358398 3220 358458
rect -960 358308 480 358398
rect 583520 351930 584960 352020
rect 580796 351870 584960 351930
rect 583520 351780 584960 351870
rect -960 345402 480 345492
rect 1534 345478 3220 345538
rect 1534 345402 1594 345478
rect -960 345342 1594 345402
rect -960 345252 480 345342
rect 580766 338602 580826 338844
rect 583520 338602 584960 338692
rect 580766 338542 584960 338602
rect 583520 338452 584960 338542
rect -960 332346 480 332436
rect 3190 332346 3250 332724
rect -960 332286 3250 332346
rect -960 332196 480 332286
rect 580766 325274 580826 325788
rect 583520 325274 584960 325364
rect 580766 325214 584960 325274
rect 583520 325124 584960 325214
rect -960 319290 480 319380
rect 3190 319290 3250 319940
rect -960 319230 3250 319290
rect -960 319140 480 319230
rect 580766 312082 580826 312732
rect 583520 312082 584960 312172
rect 580766 312022 584960 312082
rect 583520 311932 584960 312022
rect -960 306234 480 306324
rect 3190 306234 3250 307156
rect -960 306174 3250 306234
rect -960 306084 480 306174
rect 580766 299298 580826 299676
rect 580766 299238 583586 299298
rect 583526 298890 583586 299238
rect 583342 298844 583586 298890
rect 583342 298830 584960 298844
rect 583342 298754 583402 298830
rect 583520 298754 584960 298830
rect 583342 298694 584960 298754
rect 583520 298604 584960 298694
rect 1301 294402 1367 294405
rect 1301 294400 3220 294402
rect 1301 294344 1306 294400
rect 1362 294344 3220 294400
rect 1301 294342 3220 294344
rect 1301 294339 1367 294342
rect -960 293178 480 293268
rect 1301 293178 1367 293181
rect -960 293176 1367 293178
rect -960 293120 1306 293176
rect 1362 293120 1367 293176
rect -960 293118 1367 293120
rect -960 293028 480 293118
rect 1301 293115 1367 293118
rect 580766 285970 580826 286620
rect 580766 285910 583586 285970
rect 583526 285562 583586 285910
rect 583342 285516 583586 285562
rect 583342 285502 584960 285516
rect 583342 285426 583402 285502
rect 583520 285426 584960 285502
rect 583342 285366 584960 285426
rect 583520 285276 584960 285366
rect 2773 281618 2839 281621
rect 2773 281616 3220 281618
rect 2773 281560 2778 281616
rect 2834 281560 3220 281616
rect 2773 281558 3220 281560
rect 2773 281555 2839 281558
rect -960 280122 480 280212
rect 2773 280122 2839 280125
rect -960 280120 2839 280122
rect -960 280064 2778 280120
rect 2834 280064 2839 280120
rect -960 280062 2839 280064
rect -960 279972 480 280062
rect 2773 280059 2839 280062
rect 580766 272914 580826 273564
rect 580766 272854 583586 272914
rect 583526 272370 583586 272854
rect 583342 272324 583586 272370
rect 583342 272310 584960 272324
rect 583342 272234 583402 272310
rect 583520 272234 584960 272310
rect 583342 272174 584960 272234
rect 583520 272084 584960 272174
rect 1301 268834 1367 268837
rect 1301 268832 3220 268834
rect 1301 268776 1306 268832
rect 1362 268776 3220 268832
rect 1301 268774 3220 268776
rect 1301 268771 1367 268774
rect -960 267202 480 267292
rect 1301 267202 1367 267205
rect -960 267200 1367 267202
rect -960 267144 1306 267200
rect 1362 267144 1367 267200
rect -960 267142 1367 267144
rect -960 267052 480 267142
rect 1301 267139 1367 267142
rect 582373 260538 582439 260541
rect 580796 260536 582439 260538
rect 580796 260480 582378 260536
rect 582434 260480 582439 260536
rect 580796 260478 582439 260480
rect 582373 260475 582439 260478
rect 582373 258906 582439 258909
rect 583520 258906 584960 258996
rect 582373 258904 584960 258906
rect 582373 258848 582378 258904
rect 582434 258848 584960 258904
rect 582373 258846 584960 258848
rect 582373 258843 582439 258846
rect 583520 258756 584960 258846
rect 1301 256050 1367 256053
rect 1301 256048 3220 256050
rect 1301 255992 1306 256048
rect 1362 255992 3220 256048
rect 1301 255990 3220 255992
rect 1301 255987 1367 255990
rect -960 254146 480 254236
rect 1301 254146 1367 254149
rect -960 254144 1367 254146
rect -960 254088 1306 254144
rect 1362 254088 1367 254144
rect -960 254086 1367 254088
rect -960 253996 480 254086
rect 1301 254083 1367 254086
rect 580766 247074 580826 247452
rect 580901 247074 580967 247077
rect 580766 247072 580967 247074
rect 580766 247016 580906 247072
rect 580962 247016 580967 247072
rect 580766 247014 580967 247016
rect 580901 247011 580967 247014
rect 580901 245578 580967 245581
rect 583520 245578 584960 245668
rect 580901 245576 584960 245578
rect 580901 245520 580906 245576
rect 580962 245520 584960 245576
rect 580901 245518 584960 245520
rect 580901 245515 580967 245518
rect 583520 245428 584960 245518
rect 2773 243266 2839 243269
rect 2773 243264 3220 243266
rect 2773 243208 2778 243264
rect 2834 243208 3220 243264
rect 2773 243206 3220 243208
rect 2773 243203 2839 243206
rect -960 241090 480 241180
rect 2773 241090 2839 241093
rect -960 241088 2839 241090
rect -960 241032 2778 241088
rect 2834 241032 2839 241088
rect -960 241030 2839 241032
rect -960 240940 480 241030
rect 2773 241027 2839 241030
rect 582373 234426 582439 234429
rect 580796 234424 582439 234426
rect 580796 234368 582378 234424
rect 582434 234368 582439 234424
rect 580796 234366 582439 234368
rect 582373 234363 582439 234366
rect 582373 232386 582439 232389
rect 583520 232386 584960 232476
rect 582373 232384 584960 232386
rect 582373 232328 582378 232384
rect 582434 232328 584960 232384
rect 582373 232326 584960 232328
rect 582373 232323 582439 232326
rect 583520 232236 584960 232326
rect 2773 230618 2839 230621
rect 2773 230616 3220 230618
rect 2773 230560 2778 230616
rect 2834 230560 3220 230616
rect 2773 230558 3220 230560
rect 2773 230555 2839 230558
rect -960 228034 480 228124
rect 2773 228034 2839 228037
rect -960 228032 2839 228034
rect -960 227976 2778 228032
rect 2834 227976 2839 228032
rect -960 227974 2839 227976
rect -960 227884 480 227974
rect 2773 227971 2839 227974
rect 580766 220962 580826 221340
rect 580901 220962 580967 220965
rect 580766 220960 580967 220962
rect 580766 220904 580906 220960
rect 580962 220904 580967 220960
rect 580766 220902 580967 220904
rect 580901 220899 580967 220902
rect 580901 219058 580967 219061
rect 583520 219058 584960 219148
rect 580901 219056 584960 219058
rect 580901 219000 580906 219056
rect 580962 219000 584960 219056
rect 580901 218998 584960 219000
rect 580901 218995 580967 218998
rect 583520 218908 584960 218998
rect 2773 217698 2839 217701
rect 2773 217696 3220 217698
rect 2773 217640 2778 217696
rect 2834 217640 3220 217696
rect 2773 217638 3220 217640
rect 2773 217635 2839 217638
rect -960 214978 480 215068
rect 2773 214978 2839 214981
rect -960 214976 2839 214978
rect -960 214920 2778 214976
rect 2834 214920 2839 214976
rect -960 214918 2839 214920
rect -960 214828 480 214918
rect 2773 214915 2839 214918
rect 582373 208314 582439 208317
rect 580796 208312 582439 208314
rect 580796 208256 582378 208312
rect 582434 208256 582439 208312
rect 580796 208254 582439 208256
rect 582373 208251 582439 208254
rect 582373 205730 582439 205733
rect 583520 205730 584960 205820
rect 582373 205728 584960 205730
rect 582373 205672 582378 205728
rect 582434 205672 584960 205728
rect 582373 205670 584960 205672
rect 582373 205667 582439 205670
rect 583520 205580 584960 205670
rect 2773 204914 2839 204917
rect 2773 204912 3220 204914
rect 2773 204856 2778 204912
rect 2834 204856 3220 204912
rect 2773 204854 3220 204856
rect 2773 204851 2839 204854
rect -960 201922 480 202012
rect 2773 201922 2839 201925
rect -960 201920 2839 201922
rect -960 201864 2778 201920
rect 2834 201864 2839 201920
rect -960 201862 2839 201864
rect -960 201772 480 201862
rect 2773 201859 2839 201862
rect 580766 194714 580826 195228
rect 580901 194714 580967 194717
rect 580766 194712 580967 194714
rect 580766 194656 580906 194712
rect 580962 194656 580967 194712
rect 580766 194654 580967 194656
rect 580901 194651 580967 194654
rect 580901 192538 580967 192541
rect 583520 192538 584960 192628
rect 580901 192536 584960 192538
rect 580901 192480 580906 192536
rect 580962 192480 584960 192536
rect 580901 192478 584960 192480
rect 580901 192475 580967 192478
rect 583520 192388 584960 192478
rect 1301 192130 1367 192133
rect 1301 192128 3220 192130
rect 1301 192072 1306 192128
rect 1362 192072 3220 192128
rect 1301 192070 3220 192072
rect 1301 192067 1367 192070
rect -960 188866 480 188956
rect 1301 188866 1367 188869
rect -960 188864 1367 188866
rect -960 188808 1306 188864
rect 1362 188808 1367 188864
rect -960 188806 1367 188808
rect -960 188716 480 188806
rect 1301 188803 1367 188806
rect 580901 182474 580967 182477
rect 580766 182472 580967 182474
rect 580766 182416 580906 182472
rect 580962 182416 580967 182472
rect 580766 182414 580967 182416
rect 580766 182308 580826 182414
rect 580901 182411 580967 182414
rect 2773 179346 2839 179349
rect 2773 179344 3220 179346
rect 2773 179288 2778 179344
rect 2834 179288 3220 179344
rect 2773 179286 3220 179288
rect 2773 179283 2839 179286
rect 580901 179210 580967 179213
rect 583520 179210 584960 179300
rect 580901 179208 584960 179210
rect 580901 179152 580906 179208
rect 580962 179152 584960 179208
rect 580901 179150 584960 179152
rect 580901 179147 580967 179150
rect 583520 179060 584960 179150
rect -960 175946 480 176036
rect 2773 175946 2839 175949
rect -960 175944 2839 175946
rect -960 175888 2778 175944
rect 2834 175888 2839 175944
rect -960 175886 2839 175888
rect -960 175796 480 175886
rect 2773 175883 2839 175886
rect 580766 168602 580826 169116
rect 580901 168602 580967 168605
rect 580766 168600 580967 168602
rect 580766 168544 580906 168600
rect 580962 168544 580967 168600
rect 580766 168542 580967 168544
rect 580901 168539 580967 168542
rect 2773 166562 2839 166565
rect 2773 166560 3220 166562
rect 2773 166504 2778 166560
rect 2834 166504 3220 166560
rect 2773 166502 3220 166504
rect 2773 166499 2839 166502
rect 580901 165882 580967 165885
rect 583520 165882 584960 165972
rect 580901 165880 584960 165882
rect 580901 165824 580906 165880
rect 580962 165824 584960 165880
rect 580901 165822 584960 165824
rect 580901 165819 580967 165822
rect 583520 165732 584960 165822
rect -960 162890 480 162980
rect 2773 162890 2839 162893
rect -960 162888 2839 162890
rect -960 162832 2778 162888
rect 2834 162832 2839 162888
rect -960 162830 2839 162832
rect -960 162740 480 162830
rect 2773 162827 2839 162830
rect 580901 156362 580967 156365
rect 580766 156360 580967 156362
rect 580766 156304 580906 156360
rect 580962 156304 580967 156360
rect 580766 156302 580967 156304
rect 580766 156196 580826 156302
rect 580901 156299 580967 156302
rect 1301 153778 1367 153781
rect 1301 153776 3220 153778
rect 1301 153720 1306 153776
rect 1362 153720 3220 153776
rect 1301 153718 3220 153720
rect 1301 153715 1367 153718
rect 580901 152690 580967 152693
rect 583520 152690 584960 152780
rect 580901 152688 584960 152690
rect 580901 152632 580906 152688
rect 580962 152632 584960 152688
rect 580901 152630 584960 152632
rect 580901 152627 580967 152630
rect 583520 152540 584960 152630
rect -960 149834 480 149924
rect 1301 149834 1367 149837
rect -960 149832 1367 149834
rect -960 149776 1306 149832
rect 1362 149776 1367 149832
rect -960 149774 1367 149776
rect -960 149684 480 149774
rect 1301 149771 1367 149774
rect 580766 142626 580826 143004
rect 580901 142626 580967 142629
rect 580766 142624 580967 142626
rect 580766 142568 580906 142624
rect 580962 142568 580967 142624
rect 580766 142566 580967 142568
rect 580901 142563 580967 142566
rect 565 140994 631 140997
rect 565 140992 3220 140994
rect 565 140936 570 140992
rect 626 140936 3220 140992
rect 565 140934 3220 140936
rect 565 140931 631 140934
rect 580901 139362 580967 139365
rect 583520 139362 584960 139452
rect 580901 139360 584960 139362
rect 580901 139304 580906 139360
rect 580962 139304 584960 139360
rect 580901 139302 584960 139304
rect 580901 139299 580967 139302
rect 583520 139212 584960 139302
rect -960 136778 480 136868
rect 565 136778 631 136781
rect -960 136776 631 136778
rect -960 136720 570 136776
rect 626 136720 631 136776
rect -960 136718 631 136720
rect -960 136628 480 136718
rect 565 136715 631 136718
rect 580901 130250 580967 130253
rect 580766 130248 580967 130250
rect 580766 130192 580906 130248
rect 580962 130192 580967 130248
rect 580766 130190 580967 130192
rect 580766 130084 580826 130190
rect 580901 130187 580967 130190
rect 749 128210 815 128213
rect 749 128208 3220 128210
rect 749 128152 754 128208
rect 810 128152 3220 128208
rect 749 128150 3220 128152
rect 749 128147 815 128150
rect 580901 126034 580967 126037
rect 583520 126034 584960 126124
rect 580901 126032 584960 126034
rect 580901 125976 580906 126032
rect 580962 125976 584960 126032
rect 580901 125974 584960 125976
rect 580901 125971 580967 125974
rect 583520 125884 584960 125974
rect -960 123722 480 123812
rect 749 123722 815 123725
rect -960 123720 815 123722
rect -960 123664 754 123720
rect 810 123664 815 123720
rect -960 123662 815 123664
rect -960 123572 480 123662
rect 749 123659 815 123662
rect 579889 116378 579955 116381
rect 580030 116378 580090 116892
rect 579889 116376 580090 116378
rect 579889 116320 579894 116376
rect 579950 116320 580090 116376
rect 579889 116318 580090 116320
rect 579889 116315 579955 116318
rect 1301 115426 1367 115429
rect 1301 115424 3220 115426
rect 1301 115368 1306 115424
rect 1362 115368 3220 115424
rect 1301 115366 3220 115368
rect 1301 115363 1367 115366
rect 579889 112842 579955 112845
rect 583520 112842 584960 112932
rect 579889 112840 584960 112842
rect 579889 112784 579894 112840
rect 579950 112784 584960 112840
rect 579889 112782 584960 112784
rect 579889 112779 579955 112782
rect 583520 112692 584960 112782
rect -960 110666 480 110756
rect 1301 110666 1367 110669
rect -960 110664 1367 110666
rect -960 110608 1306 110664
rect 1362 110608 1367 110664
rect -960 110606 1367 110608
rect -960 110516 480 110606
rect 1301 110603 1367 110606
rect 580766 103594 580826 103836
rect 580901 103594 580967 103597
rect 580766 103592 580967 103594
rect 580766 103536 580906 103592
rect 580962 103536 580967 103592
rect 580766 103534 580967 103536
rect 580901 103531 580967 103534
rect 1577 102642 1643 102645
rect 1577 102640 3220 102642
rect 1577 102584 1582 102640
rect 1638 102584 3220 102640
rect 1577 102582 3220 102584
rect 1577 102579 1643 102582
rect 580901 99514 580967 99517
rect 583520 99514 584960 99604
rect 580901 99512 584960 99514
rect 580901 99456 580906 99512
rect 580962 99456 584960 99512
rect 580901 99454 584960 99456
rect 580901 99451 580967 99454
rect 583520 99364 584960 99454
rect -960 97610 480 97700
rect 1577 97610 1643 97613
rect -960 97608 1643 97610
rect -960 97552 1582 97608
rect 1638 97552 1643 97608
rect -960 97550 1643 97552
rect -960 97460 480 97550
rect 1577 97547 1643 97550
rect 580766 90266 580826 90780
rect 580901 90266 580967 90269
rect 580766 90264 580967 90266
rect 580766 90208 580906 90264
rect 580962 90208 580967 90264
rect 580766 90206 580967 90208
rect 580901 90203 580967 90206
rect 1577 89858 1643 89861
rect 1577 89856 3220 89858
rect 1577 89800 1582 89856
rect 1638 89800 3220 89856
rect 1577 89798 3220 89800
rect 1577 89795 1643 89798
rect 580901 86186 580967 86189
rect 583520 86186 584960 86276
rect 580901 86184 584960 86186
rect 580901 86128 580906 86184
rect 580962 86128 584960 86184
rect 580901 86126 584960 86128
rect 580901 86123 580967 86126
rect 583520 86036 584960 86126
rect -960 84690 480 84780
rect 1577 84690 1643 84693
rect -960 84688 1643 84690
rect -960 84632 1582 84688
rect 1638 84632 1643 84688
rect -960 84630 1643 84632
rect -960 84540 480 84630
rect 1577 84627 1643 84630
rect 579889 77346 579955 77349
rect 580030 77346 580090 77724
rect 579889 77344 580090 77346
rect 579889 77288 579894 77344
rect 579950 77288 580090 77344
rect 579889 77286 580090 77288
rect 579889 77283 579955 77286
rect 1577 77074 1643 77077
rect 1577 77072 3220 77074
rect 1577 77016 1582 77072
rect 1638 77016 3220 77072
rect 1577 77014 3220 77016
rect 1577 77011 1643 77014
rect 579889 72994 579955 72997
rect 583520 72994 584960 73084
rect 579889 72992 584960 72994
rect 579889 72936 579894 72992
rect 579950 72936 584960 72992
rect 579889 72934 584960 72936
rect 579889 72931 579955 72934
rect 583520 72844 584960 72934
rect -960 71634 480 71724
rect 1577 71634 1643 71637
rect -960 71632 1643 71634
rect -960 71576 1582 71632
rect 1638 71576 1643 71632
rect -960 71574 1643 71576
rect -960 71484 480 71574
rect 1577 71571 1643 71574
rect 1485 64290 1551 64293
rect 1485 64288 3220 64290
rect 1485 64232 1490 64288
rect 1546 64232 3220 64288
rect 1485 64230 3220 64232
rect 1485 64227 1551 64230
rect 580766 64154 580826 64668
rect 580901 64154 580967 64157
rect 580766 64152 580967 64154
rect 580766 64096 580906 64152
rect 580962 64096 580967 64152
rect 580766 64094 580967 64096
rect 580901 64091 580967 64094
rect 580901 59666 580967 59669
rect 583520 59666 584960 59756
rect 580901 59664 584960 59666
rect 580901 59608 580906 59664
rect 580962 59608 584960 59664
rect 580901 59606 584960 59608
rect 580901 59603 580967 59606
rect 583520 59516 584960 59606
rect -960 58578 480 58668
rect 1485 58578 1551 58581
rect -960 58576 1551 58578
rect -960 58520 1490 58576
rect 1546 58520 1551 58576
rect -960 58518 1551 58520
rect -960 58428 480 58518
rect 1485 58515 1551 58518
rect 2037 51506 2103 51509
rect 2037 51504 3220 51506
rect 2037 51448 2042 51504
rect 2098 51448 3220 51504
rect 2037 51446 3220 51448
rect 2037 51443 2103 51446
rect 580766 51098 580826 51612
rect 580901 51098 580967 51101
rect 580766 51096 580967 51098
rect 580766 51040 580906 51096
rect 580962 51040 580967 51096
rect 580766 51038 580967 51040
rect 580901 51035 580967 51038
rect 580901 46338 580967 46341
rect 583520 46338 584960 46428
rect 580901 46336 584960 46338
rect 580901 46280 580906 46336
rect 580962 46280 584960 46336
rect 580901 46278 584960 46280
rect 580901 46275 580967 46278
rect 583520 46188 584960 46278
rect -960 45522 480 45612
rect 2037 45522 2103 45525
rect -960 45520 2103 45522
rect -960 45464 2042 45520
rect 2098 45464 2103 45520
rect -960 45462 2103 45464
rect -960 45372 480 45462
rect 2037 45459 2103 45462
rect 2037 38722 2103 38725
rect 2037 38720 3220 38722
rect 2037 38664 2042 38720
rect 2098 38664 3220 38720
rect 2037 38662 3220 38664
rect 2037 38659 2103 38662
rect 580766 38042 580826 38556
rect 580901 38042 580967 38045
rect 580766 38040 580967 38042
rect 580766 37984 580906 38040
rect 580962 37984 580967 38040
rect 580766 37982 580967 37984
rect 580901 37979 580967 37982
rect 580901 33146 580967 33149
rect 583520 33146 584960 33236
rect 580901 33144 584960 33146
rect 580901 33088 580906 33144
rect 580962 33088 584960 33144
rect 580901 33086 584960 33088
rect 580901 33083 580967 33086
rect 583520 32996 584960 33086
rect -960 32466 480 32556
rect 2037 32466 2103 32469
rect -960 32464 2103 32466
rect -960 32408 2042 32464
rect 2098 32408 2103 32464
rect -960 32406 2103 32408
rect -960 32316 480 32406
rect 2037 32403 2103 32406
rect 1485 25938 1551 25941
rect 1485 25936 3220 25938
rect 1485 25880 1490 25936
rect 1546 25880 3220 25936
rect 1485 25878 3220 25880
rect 1485 25875 1551 25878
rect 580766 24986 580826 25500
rect 580901 24986 580967 24989
rect 580766 24984 580967 24986
rect 580766 24928 580906 24984
rect 580962 24928 580967 24984
rect 580766 24926 580967 24928
rect 580901 24923 580967 24926
rect 580901 19818 580967 19821
rect 583520 19818 584960 19908
rect 580901 19816 584960 19818
rect 580901 19760 580906 19816
rect 580962 19760 584960 19816
rect 580901 19758 584960 19760
rect 580901 19755 580967 19758
rect 583520 19668 584960 19758
rect -960 19410 480 19500
rect 1485 19410 1551 19413
rect -960 19408 1551 19410
rect -960 19352 1490 19408
rect 1546 19352 1551 19408
rect -960 19350 1551 19352
rect -960 19260 480 19350
rect 1485 19347 1551 19350
rect 2037 13154 2103 13157
rect 2037 13152 3220 13154
rect 2037 13096 2042 13152
rect 2098 13096 3220 13152
rect 2037 13094 3220 13096
rect 2037 13091 2103 13094
rect 579889 12746 579955 12749
rect 579889 12744 580090 12746
rect 579889 12688 579894 12744
rect 579950 12688 580090 12744
rect 579889 12686 580090 12688
rect 579889 12683 579955 12686
rect 580030 12580 580090 12686
rect 579889 6626 579955 6629
rect 583520 6626 584960 6716
rect 579889 6624 584960 6626
rect -960 6490 480 6580
rect 579889 6568 579894 6624
rect 579950 6568 584960 6624
rect 579889 6566 584960 6568
rect 579889 6563 579955 6566
rect 2037 6490 2103 6493
rect -960 6488 2103 6490
rect -960 6432 2042 6488
rect 2098 6432 2103 6488
rect 583520 6476 584960 6566
rect -960 6430 2103 6432
rect -960 6340 480 6430
rect 2037 6427 2103 6430
rect 70209 3906 70275 3909
rect 73613 3906 73679 3909
rect 70209 3904 73679 3906
rect 70209 3848 70214 3904
rect 70270 3848 73618 3904
rect 73674 3848 73679 3904
rect 70209 3846 73679 3848
rect 70209 3843 70275 3846
rect 73613 3843 73679 3846
rect 28901 642 28967 645
rect 46289 642 46355 645
rect 28901 640 46355 642
rect 28901 584 28906 640
rect 28962 584 46294 640
rect 46350 584 46355 640
rect 28901 582 46355 584
rect 28901 579 28967 582
rect 46289 579 46355 582
rect 12157 506 12223 509
rect 30833 506 30899 509
rect 12157 504 30899 506
rect 12157 448 12162 504
rect 12218 448 30838 504
rect 30894 448 30899 504
rect 12157 446 30899 448
rect 12157 443 12223 446
rect 30833 443 30899 446
rect 5441 370 5507 373
rect 23933 370 23999 373
rect 5441 368 23999 370
rect 5441 312 5446 368
rect 5502 312 23938 368
rect 23994 312 23999 368
rect 5441 310 23999 312
rect 5441 307 5507 310
rect 23933 307 23999 310
rect 25681 370 25747 373
rect 42701 370 42767 373
rect 25681 368 42767 370
rect 25681 312 25686 368
rect 25742 312 42706 368
rect 42762 312 42767 368
rect 25681 310 42767 312
rect 25681 307 25747 310
rect 42701 307 42767 310
rect 13721 234 13787 237
rect 31937 234 32003 237
rect 13721 232 32003 234
rect 13721 176 13726 232
rect 13782 176 31942 232
rect 31998 176 32003 232
rect 13721 174 32003 176
rect 13721 171 13787 174
rect 31937 171 32003 174
rect 36997 234 37063 237
rect 54017 234 54083 237
rect 36997 232 54083 234
rect 36997 176 37002 232
rect 37058 176 54022 232
rect 54078 176 54083 232
rect 36997 174 54083 176
rect 36997 171 37063 174
rect 54017 171 54083 174
rect 6269 98 6335 101
rect 25037 98 25103 101
rect 6269 96 25103 98
rect 6269 40 6274 96
rect 6330 40 25042 96
rect 25098 40 25103 96
rect 6269 38 25103 40
rect 6269 35 6335 38
rect 25037 35 25103 38
rect 46841 98 46907 101
rect 62849 98 62915 101
rect 46841 96 62915 98
rect 46841 40 46846 96
rect 46902 40 62854 96
rect 62910 40 62915 96
rect 46841 38 62915 40
rect 46841 35 46907 38
rect 62849 35 62915 38
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 -7066 -8106 711002
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 -6106 -7146 710042
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 -5146 -6186 709082
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 -4186 -5226 708122
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 -3226 -4266 707162
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 -2266 -3306 706202
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 694354 -2346 705242
rect 582294 705798 582914 711590
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 582294 705562 582326 705798
rect 582562 705562 582646 705798
rect 582882 705562 582914 705798
rect 582294 705478 582914 705562
rect 582294 705242 582326 705478
rect 582562 705242 582646 705478
rect 582882 705242 582914 705478
rect -2966 694118 -2934 694354
rect -2698 694118 -2614 694354
rect -2378 694118 -2346 694354
rect -2966 694034 -2346 694118
rect -2966 693798 -2934 694034
rect -2698 693798 -2614 694034
rect -2378 693798 -2346 694034
rect -2966 658354 -2346 693798
rect -2966 658118 -2934 658354
rect -2698 658118 -2614 658354
rect -2378 658118 -2346 658354
rect -2966 658034 -2346 658118
rect -2966 657798 -2934 658034
rect -2698 657798 -2614 658034
rect -2378 657798 -2346 658034
rect -2966 622354 -2346 657798
rect -2966 622118 -2934 622354
rect -2698 622118 -2614 622354
rect -2378 622118 -2346 622354
rect -2966 622034 -2346 622118
rect -2966 621798 -2934 622034
rect -2698 621798 -2614 622034
rect -2378 621798 -2346 622034
rect -2966 586354 -2346 621798
rect -2966 586118 -2934 586354
rect -2698 586118 -2614 586354
rect -2378 586118 -2346 586354
rect -2966 586034 -2346 586118
rect -2966 585798 -2934 586034
rect -2698 585798 -2614 586034
rect -2378 585798 -2346 586034
rect -2966 550354 -2346 585798
rect -2966 550118 -2934 550354
rect -2698 550118 -2614 550354
rect -2378 550118 -2346 550354
rect -2966 550034 -2346 550118
rect -2966 549798 -2934 550034
rect -2698 549798 -2614 550034
rect -2378 549798 -2346 550034
rect -2966 514354 -2346 549798
rect -2966 514118 -2934 514354
rect -2698 514118 -2614 514354
rect -2378 514118 -2346 514354
rect -2966 514034 -2346 514118
rect -2966 513798 -2934 514034
rect -2698 513798 -2614 514034
rect -2378 513798 -2346 514034
rect -2966 478354 -2346 513798
rect -2966 478118 -2934 478354
rect -2698 478118 -2614 478354
rect -2378 478118 -2346 478354
rect -2966 478034 -2346 478118
rect -2966 477798 -2934 478034
rect -2698 477798 -2614 478034
rect -2378 477798 -2346 478034
rect -2966 442354 -2346 477798
rect -2966 442118 -2934 442354
rect -2698 442118 -2614 442354
rect -2378 442118 -2346 442354
rect -2966 442034 -2346 442118
rect -2966 441798 -2934 442034
rect -2698 441798 -2614 442034
rect -2378 441798 -2346 442034
rect -2966 406354 -2346 441798
rect -2966 406118 -2934 406354
rect -2698 406118 -2614 406354
rect -2378 406118 -2346 406354
rect -2966 406034 -2346 406118
rect -2966 405798 -2934 406034
rect -2698 405798 -2614 406034
rect -2378 405798 -2346 406034
rect -2966 370354 -2346 405798
rect -2966 370118 -2934 370354
rect -2698 370118 -2614 370354
rect -2378 370118 -2346 370354
rect -2966 370034 -2346 370118
rect -2966 369798 -2934 370034
rect -2698 369798 -2614 370034
rect -2378 369798 -2346 370034
rect -2966 334354 -2346 369798
rect -2966 334118 -2934 334354
rect -2698 334118 -2614 334354
rect -2378 334118 -2346 334354
rect -2966 334034 -2346 334118
rect -2966 333798 -2934 334034
rect -2698 333798 -2614 334034
rect -2378 333798 -2346 334034
rect -2966 298354 -2346 333798
rect -2966 298118 -2934 298354
rect -2698 298118 -2614 298354
rect -2378 298118 -2346 298354
rect -2966 298034 -2346 298118
rect -2966 297798 -2934 298034
rect -2698 297798 -2614 298034
rect -2378 297798 -2346 298034
rect -2966 262354 -2346 297798
rect -2966 262118 -2934 262354
rect -2698 262118 -2614 262354
rect -2378 262118 -2346 262354
rect -2966 262034 -2346 262118
rect -2966 261798 -2934 262034
rect -2698 261798 -2614 262034
rect -2378 261798 -2346 262034
rect -2966 226354 -2346 261798
rect -2966 226118 -2934 226354
rect -2698 226118 -2614 226354
rect -2378 226118 -2346 226354
rect -2966 226034 -2346 226118
rect -2966 225798 -2934 226034
rect -2698 225798 -2614 226034
rect -2378 225798 -2346 226034
rect -2966 190354 -2346 225798
rect -2966 190118 -2934 190354
rect -2698 190118 -2614 190354
rect -2378 190118 -2346 190354
rect -2966 190034 -2346 190118
rect -2966 189798 -2934 190034
rect -2698 189798 -2614 190034
rect -2378 189798 -2346 190034
rect -2966 154354 -2346 189798
rect -2966 154118 -2934 154354
rect -2698 154118 -2614 154354
rect -2378 154118 -2346 154354
rect -2966 154034 -2346 154118
rect -2966 153798 -2934 154034
rect -2698 153798 -2614 154034
rect -2378 153798 -2346 154034
rect -2966 118354 -2346 153798
rect -2966 118118 -2934 118354
rect -2698 118118 -2614 118354
rect -2378 118118 -2346 118354
rect -2966 118034 -2346 118118
rect -2966 117798 -2934 118034
rect -2698 117798 -2614 118034
rect -2378 117798 -2346 118034
rect -2966 82354 -2346 117798
rect -2966 82118 -2934 82354
rect -2698 82118 -2614 82354
rect -2378 82118 -2346 82354
rect -2966 82034 -2346 82118
rect -2966 81798 -2934 82034
rect -2698 81798 -2614 82034
rect -2378 81798 -2346 82034
rect -2966 46354 -2346 81798
rect -2966 46118 -2934 46354
rect -2698 46118 -2614 46354
rect -2378 46118 -2346 46354
rect -2966 46034 -2346 46118
rect -2966 45798 -2934 46034
rect -2698 45798 -2614 46034
rect -2378 45798 -2346 46034
rect -2966 10354 -2346 45798
rect -2966 10118 -2934 10354
rect -2698 10118 -2614 10354
rect -2378 10118 -2346 10354
rect -2966 10034 -2346 10118
rect -2966 9798 -2934 10034
rect -2698 9798 -2614 10034
rect -2378 9798 -2346 10034
rect -2966 -1306 -2346 9798
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 689854 -1386 704282
rect 582294 694354 582914 705242
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 23794 694118 23826 694354
rect 24062 694118 24146 694354
rect 24382 694118 24414 694354
rect 23794 694034 24414 694118
rect 23794 693798 23826 694034
rect 24062 693798 24146 694034
rect 24382 693798 24414 694034
rect 59794 694118 59826 694354
rect 60062 694118 60146 694354
rect 60382 694118 60414 694354
rect 59794 694034 60414 694118
rect 59794 693798 59826 694034
rect 60062 693798 60146 694034
rect 60382 693798 60414 694034
rect 95794 694118 95826 694354
rect 96062 694118 96146 694354
rect 96382 694118 96414 694354
rect 95794 694034 96414 694118
rect 95794 693798 95826 694034
rect 96062 693798 96146 694034
rect 96382 693798 96414 694034
rect 131794 694118 131826 694354
rect 132062 694118 132146 694354
rect 132382 694118 132414 694354
rect 131794 694034 132414 694118
rect 131794 693798 131826 694034
rect 132062 693798 132146 694034
rect 132382 693798 132414 694034
rect 167794 694118 167826 694354
rect 168062 694118 168146 694354
rect 168382 694118 168414 694354
rect 167794 694034 168414 694118
rect 167794 693798 167826 694034
rect 168062 693798 168146 694034
rect 168382 693798 168414 694034
rect 203794 694118 203826 694354
rect 204062 694118 204146 694354
rect 204382 694118 204414 694354
rect 203794 694034 204414 694118
rect 203794 693798 203826 694034
rect 204062 693798 204146 694034
rect 204382 693798 204414 694034
rect 239794 694118 239826 694354
rect 240062 694118 240146 694354
rect 240382 694118 240414 694354
rect 239794 694034 240414 694118
rect 239794 693798 239826 694034
rect 240062 693798 240146 694034
rect 240382 693798 240414 694034
rect 275794 694118 275826 694354
rect 276062 694118 276146 694354
rect 276382 694118 276414 694354
rect 275794 694034 276414 694118
rect 275794 693798 275826 694034
rect 276062 693798 276146 694034
rect 276382 693798 276414 694034
rect 311794 694118 311826 694354
rect 312062 694118 312146 694354
rect 312382 694118 312414 694354
rect 311794 694034 312414 694118
rect 311794 693798 311826 694034
rect 312062 693798 312146 694034
rect 312382 693798 312414 694034
rect 347794 694118 347826 694354
rect 348062 694118 348146 694354
rect 348382 694118 348414 694354
rect 347794 694034 348414 694118
rect 347794 693798 347826 694034
rect 348062 693798 348146 694034
rect 348382 693798 348414 694034
rect 383794 694118 383826 694354
rect 384062 694118 384146 694354
rect 384382 694118 384414 694354
rect 383794 694034 384414 694118
rect 383794 693798 383826 694034
rect 384062 693798 384146 694034
rect 384382 693798 384414 694034
rect 419794 694118 419826 694354
rect 420062 694118 420146 694354
rect 420382 694118 420414 694354
rect 419794 694034 420414 694118
rect 419794 693798 419826 694034
rect 420062 693798 420146 694034
rect 420382 693798 420414 694034
rect 455794 694118 455826 694354
rect 456062 694118 456146 694354
rect 456382 694118 456414 694354
rect 455794 694034 456414 694118
rect 455794 693798 455826 694034
rect 456062 693798 456146 694034
rect 456382 693798 456414 694034
rect 491794 694118 491826 694354
rect 492062 694118 492146 694354
rect 492382 694118 492414 694354
rect 491794 694034 492414 694118
rect 491794 693798 491826 694034
rect 492062 693798 492146 694034
rect 492382 693798 492414 694034
rect 527794 694118 527826 694354
rect 528062 694118 528146 694354
rect 528382 694118 528414 694354
rect 527794 694034 528414 694118
rect 527794 693798 527826 694034
rect 528062 693798 528146 694034
rect 528382 693798 528414 694034
rect 563794 694118 563826 694354
rect 564062 694118 564146 694354
rect 564382 694118 564414 694354
rect 563794 694034 564414 694118
rect 563794 693798 563826 694034
rect 564062 693798 564146 694034
rect 564382 693798 564414 694034
rect 582294 694118 582326 694354
rect 582562 694118 582646 694354
rect 582882 694118 582914 694354
rect 582294 694034 582914 694118
rect 582294 693798 582326 694034
rect 582562 693798 582646 694034
rect 582882 693798 582914 694034
rect -2006 689618 -1974 689854
rect -1738 689618 -1654 689854
rect -1418 689618 -1386 689854
rect -2006 689534 -1386 689618
rect -2006 689298 -1974 689534
rect -1738 689298 -1654 689534
rect -1418 689298 -1386 689534
rect 5794 689618 5826 689854
rect 6062 689618 6146 689854
rect 6382 689618 6414 689854
rect 5794 689534 6414 689618
rect 5794 689298 5826 689534
rect 6062 689298 6146 689534
rect 6382 689298 6414 689534
rect 41794 689618 41826 689854
rect 42062 689618 42146 689854
rect 42382 689618 42414 689854
rect 41794 689534 42414 689618
rect 41794 689298 41826 689534
rect 42062 689298 42146 689534
rect 42382 689298 42414 689534
rect 77794 689618 77826 689854
rect 78062 689618 78146 689854
rect 78382 689618 78414 689854
rect 77794 689534 78414 689618
rect 77794 689298 77826 689534
rect 78062 689298 78146 689534
rect 78382 689298 78414 689534
rect 113794 689618 113826 689854
rect 114062 689618 114146 689854
rect 114382 689618 114414 689854
rect 113794 689534 114414 689618
rect 113794 689298 113826 689534
rect 114062 689298 114146 689534
rect 114382 689298 114414 689534
rect 149794 689618 149826 689854
rect 150062 689618 150146 689854
rect 150382 689618 150414 689854
rect 149794 689534 150414 689618
rect 149794 689298 149826 689534
rect 150062 689298 150146 689534
rect 150382 689298 150414 689534
rect 185794 689618 185826 689854
rect 186062 689618 186146 689854
rect 186382 689618 186414 689854
rect 185794 689534 186414 689618
rect 185794 689298 185826 689534
rect 186062 689298 186146 689534
rect 186382 689298 186414 689534
rect 221794 689618 221826 689854
rect 222062 689618 222146 689854
rect 222382 689618 222414 689854
rect 221794 689534 222414 689618
rect 221794 689298 221826 689534
rect 222062 689298 222146 689534
rect 222382 689298 222414 689534
rect 257794 689618 257826 689854
rect 258062 689618 258146 689854
rect 258382 689618 258414 689854
rect 257794 689534 258414 689618
rect 257794 689298 257826 689534
rect 258062 689298 258146 689534
rect 258382 689298 258414 689534
rect 293794 689618 293826 689854
rect 294062 689618 294146 689854
rect 294382 689618 294414 689854
rect 293794 689534 294414 689618
rect 293794 689298 293826 689534
rect 294062 689298 294146 689534
rect 294382 689298 294414 689534
rect 329794 689618 329826 689854
rect 330062 689618 330146 689854
rect 330382 689618 330414 689854
rect 329794 689534 330414 689618
rect 329794 689298 329826 689534
rect 330062 689298 330146 689534
rect 330382 689298 330414 689534
rect 365794 689618 365826 689854
rect 366062 689618 366146 689854
rect 366382 689618 366414 689854
rect 365794 689534 366414 689618
rect 365794 689298 365826 689534
rect 366062 689298 366146 689534
rect 366382 689298 366414 689534
rect 401794 689618 401826 689854
rect 402062 689618 402146 689854
rect 402382 689618 402414 689854
rect 401794 689534 402414 689618
rect 401794 689298 401826 689534
rect 402062 689298 402146 689534
rect 402382 689298 402414 689534
rect 437794 689618 437826 689854
rect 438062 689618 438146 689854
rect 438382 689618 438414 689854
rect 437794 689534 438414 689618
rect 437794 689298 437826 689534
rect 438062 689298 438146 689534
rect 438382 689298 438414 689534
rect 473794 689618 473826 689854
rect 474062 689618 474146 689854
rect 474382 689618 474414 689854
rect 473794 689534 474414 689618
rect 473794 689298 473826 689534
rect 474062 689298 474146 689534
rect 474382 689298 474414 689534
rect 509794 689618 509826 689854
rect 510062 689618 510146 689854
rect 510382 689618 510414 689854
rect 509794 689534 510414 689618
rect 509794 689298 509826 689534
rect 510062 689298 510146 689534
rect 510382 689298 510414 689534
rect 545794 689618 545826 689854
rect 546062 689618 546146 689854
rect 546382 689618 546414 689854
rect 545794 689534 546414 689618
rect 545794 689298 545826 689534
rect 546062 689298 546146 689534
rect 546382 689298 546414 689534
rect -2006 653854 -1386 689298
rect 582294 658354 582914 693798
rect 13166 658118 13198 658354
rect 13434 658118 13518 658354
rect 13754 658118 13786 658354
rect 13166 658034 13786 658118
rect 13166 657798 13198 658034
rect 13434 657798 13518 658034
rect 13754 657798 13786 658034
rect 167794 658118 167826 658354
rect 168062 658118 168146 658354
rect 168382 658118 168414 658354
rect 167794 658034 168414 658118
rect 167794 657798 167826 658034
rect 168062 657798 168146 658034
rect 168382 657798 168414 658034
rect 291558 658118 291590 658354
rect 291826 658118 291910 658354
rect 292146 658118 292178 658354
rect 291558 658034 292178 658118
rect 291558 657798 291590 658034
rect 291826 657798 291910 658034
rect 292146 657798 292178 658034
rect 419794 658118 419826 658354
rect 420062 658118 420146 658354
rect 420382 658118 420414 658354
rect 419794 658034 420414 658118
rect 419794 657798 419826 658034
rect 420062 657798 420146 658034
rect 420382 657798 420414 658034
rect 563794 658118 563826 658354
rect 564062 658118 564146 658354
rect 564382 658118 564414 658354
rect 563794 658034 564414 658118
rect 563794 657798 563826 658034
rect 564062 657798 564146 658034
rect 564382 657798 564414 658034
rect 582294 658118 582326 658354
rect 582562 658118 582646 658354
rect 582882 658118 582914 658354
rect 582294 658034 582914 658118
rect 582294 657798 582326 658034
rect 582562 657798 582646 658034
rect 582882 657798 582914 658034
rect -2006 653618 -1974 653854
rect -1738 653618 -1654 653854
rect -1418 653618 -1386 653854
rect -2006 653534 -1386 653618
rect -2006 653298 -1974 653534
rect -1738 653298 -1654 653534
rect -1418 653298 -1386 653534
rect 5794 653618 5826 653854
rect 6062 653618 6146 653854
rect 6382 653618 6414 653854
rect 5794 653534 6414 653618
rect 5794 653298 5826 653534
rect 6062 653298 6146 653534
rect 6382 653298 6414 653534
rect 173062 653618 173094 653854
rect 173330 653618 173414 653854
rect 173650 653618 173682 653854
rect 173062 653534 173682 653618
rect 173062 653298 173094 653534
rect 173330 653298 173414 653534
rect 173650 653298 173682 653534
rect 293794 653618 293826 653854
rect 294062 653618 294146 653854
rect 294382 653618 294414 653854
rect 293794 653534 294414 653618
rect 293794 653298 293826 653534
rect 294062 653298 294146 653534
rect 294382 653298 294414 653534
rect 401794 653618 401826 653854
rect 402062 653618 402146 653854
rect 402382 653618 402414 653854
rect 401794 653534 402414 653618
rect 401794 653298 401826 653534
rect 402062 653298 402146 653534
rect 402382 653298 402414 653534
rect 570318 653618 570350 653854
rect 570586 653618 570670 653854
rect 570906 653618 570938 653854
rect 570318 653534 570938 653618
rect 570318 653298 570350 653534
rect 570586 653298 570670 653534
rect 570906 653298 570938 653534
rect -2006 617854 -1386 653298
rect 582294 622354 582914 657798
rect 13166 622118 13198 622354
rect 13434 622118 13518 622354
rect 13754 622118 13786 622354
rect 13166 622034 13786 622118
rect 13166 621798 13198 622034
rect 13434 621798 13518 622034
rect 13754 621798 13786 622034
rect 167794 622118 167826 622354
rect 168062 622118 168146 622354
rect 168382 622118 168414 622354
rect 167794 622034 168414 622118
rect 167794 621798 167826 622034
rect 168062 621798 168146 622034
rect 168382 621798 168414 622034
rect 291558 622118 291590 622354
rect 291826 622118 291910 622354
rect 292146 622118 292178 622354
rect 291558 622034 292178 622118
rect 291558 621798 291590 622034
rect 291826 621798 291910 622034
rect 292146 621798 292178 622034
rect 419794 622118 419826 622354
rect 420062 622118 420146 622354
rect 420382 622118 420414 622354
rect 419794 622034 420414 622118
rect 419794 621798 419826 622034
rect 420062 621798 420146 622034
rect 420382 621798 420414 622034
rect 563794 622118 563826 622354
rect 564062 622118 564146 622354
rect 564382 622118 564414 622354
rect 563794 622034 564414 622118
rect 563794 621798 563826 622034
rect 564062 621798 564146 622034
rect 564382 621798 564414 622034
rect 582294 622118 582326 622354
rect 582562 622118 582646 622354
rect 582882 622118 582914 622354
rect 582294 622034 582914 622118
rect 582294 621798 582326 622034
rect 582562 621798 582646 622034
rect 582882 621798 582914 622034
rect -2006 617618 -1974 617854
rect -1738 617618 -1654 617854
rect -1418 617618 -1386 617854
rect -2006 617534 -1386 617618
rect -2006 617298 -1974 617534
rect -1738 617298 -1654 617534
rect -1418 617298 -1386 617534
rect 5794 617618 5826 617854
rect 6062 617618 6146 617854
rect 6382 617618 6414 617854
rect 5794 617534 6414 617618
rect 5794 617298 5826 617534
rect 6062 617298 6146 617534
rect 6382 617298 6414 617534
rect 173062 617618 173094 617854
rect 173330 617618 173414 617854
rect 173650 617618 173682 617854
rect 173062 617534 173682 617618
rect 173062 617298 173094 617534
rect 173330 617298 173414 617534
rect 173650 617298 173682 617534
rect 293794 617618 293826 617854
rect 294062 617618 294146 617854
rect 294382 617618 294414 617854
rect 293794 617534 294414 617618
rect 293794 617298 293826 617534
rect 294062 617298 294146 617534
rect 294382 617298 294414 617534
rect 401794 617618 401826 617854
rect 402062 617618 402146 617854
rect 402382 617618 402414 617854
rect 401794 617534 402414 617618
rect 401794 617298 401826 617534
rect 402062 617298 402146 617534
rect 402382 617298 402414 617534
rect 570318 617618 570350 617854
rect 570586 617618 570670 617854
rect 570906 617618 570938 617854
rect 570318 617534 570938 617618
rect 570318 617298 570350 617534
rect 570586 617298 570670 617534
rect 570906 617298 570938 617534
rect -2006 581854 -1386 617298
rect 582294 586354 582914 621798
rect 23794 586118 23826 586354
rect 24062 586118 24146 586354
rect 24382 586118 24414 586354
rect 23794 586034 24414 586118
rect 23794 585798 23826 586034
rect 24062 585798 24146 586034
rect 24382 585798 24414 586034
rect 59794 586118 59826 586354
rect 60062 586118 60146 586354
rect 60382 586118 60414 586354
rect 59794 586034 60414 586118
rect 59794 585798 59826 586034
rect 60062 585798 60146 586034
rect 60382 585798 60414 586034
rect 95794 586118 95826 586354
rect 96062 586118 96146 586354
rect 96382 586118 96414 586354
rect 95794 586034 96414 586118
rect 95794 585798 95826 586034
rect 96062 585798 96146 586034
rect 96382 585798 96414 586034
rect 131794 586118 131826 586354
rect 132062 586118 132146 586354
rect 132382 586118 132414 586354
rect 131794 586034 132414 586118
rect 131794 585798 131826 586034
rect 132062 585798 132146 586034
rect 132382 585798 132414 586034
rect 167794 586118 167826 586354
rect 168062 586118 168146 586354
rect 168382 586118 168414 586354
rect 167794 586034 168414 586118
rect 167794 585798 167826 586034
rect 168062 585798 168146 586034
rect 168382 585798 168414 586034
rect 203794 586118 203826 586354
rect 204062 586118 204146 586354
rect 204382 586118 204414 586354
rect 203794 586034 204414 586118
rect 203794 585798 203826 586034
rect 204062 585798 204146 586034
rect 204382 585798 204414 586034
rect 239794 586118 239826 586354
rect 240062 586118 240146 586354
rect 240382 586118 240414 586354
rect 239794 586034 240414 586118
rect 239794 585798 239826 586034
rect 240062 585798 240146 586034
rect 240382 585798 240414 586034
rect 275794 586118 275826 586354
rect 276062 586118 276146 586354
rect 276382 586118 276414 586354
rect 275794 586034 276414 586118
rect 275794 585798 275826 586034
rect 276062 585798 276146 586034
rect 276382 585798 276414 586034
rect 311794 586118 311826 586354
rect 312062 586118 312146 586354
rect 312382 586118 312414 586354
rect 311794 586034 312414 586118
rect 311794 585798 311826 586034
rect 312062 585798 312146 586034
rect 312382 585798 312414 586034
rect 347794 586118 347826 586354
rect 348062 586118 348146 586354
rect 348382 586118 348414 586354
rect 347794 586034 348414 586118
rect 347794 585798 347826 586034
rect 348062 585798 348146 586034
rect 348382 585798 348414 586034
rect 383794 586118 383826 586354
rect 384062 586118 384146 586354
rect 384382 586118 384414 586354
rect 383794 586034 384414 586118
rect 383794 585798 383826 586034
rect 384062 585798 384146 586034
rect 384382 585798 384414 586034
rect 419794 586118 419826 586354
rect 420062 586118 420146 586354
rect 420382 586118 420414 586354
rect 419794 586034 420414 586118
rect 419794 585798 419826 586034
rect 420062 585798 420146 586034
rect 420382 585798 420414 586034
rect 455794 586118 455826 586354
rect 456062 586118 456146 586354
rect 456382 586118 456414 586354
rect 455794 586034 456414 586118
rect 455794 585798 455826 586034
rect 456062 585798 456146 586034
rect 456382 585798 456414 586034
rect 491794 586118 491826 586354
rect 492062 586118 492146 586354
rect 492382 586118 492414 586354
rect 491794 586034 492414 586118
rect 491794 585798 491826 586034
rect 492062 585798 492146 586034
rect 492382 585798 492414 586034
rect 527794 586118 527826 586354
rect 528062 586118 528146 586354
rect 528382 586118 528414 586354
rect 527794 586034 528414 586118
rect 527794 585798 527826 586034
rect 528062 585798 528146 586034
rect 528382 585798 528414 586034
rect 563794 586118 563826 586354
rect 564062 586118 564146 586354
rect 564382 586118 564414 586354
rect 563794 586034 564414 586118
rect 563794 585798 563826 586034
rect 564062 585798 564146 586034
rect 564382 585798 564414 586034
rect 582294 586118 582326 586354
rect 582562 586118 582646 586354
rect 582882 586118 582914 586354
rect 582294 586034 582914 586118
rect 582294 585798 582326 586034
rect 582562 585798 582646 586034
rect 582882 585798 582914 586034
rect -2006 581618 -1974 581854
rect -1738 581618 -1654 581854
rect -1418 581618 -1386 581854
rect -2006 581534 -1386 581618
rect -2006 581298 -1974 581534
rect -1738 581298 -1654 581534
rect -1418 581298 -1386 581534
rect 5794 581618 5826 581854
rect 6062 581618 6146 581854
rect 6382 581618 6414 581854
rect 5794 581534 6414 581618
rect 5794 581298 5826 581534
rect 6062 581298 6146 581534
rect 6382 581298 6414 581534
rect 41794 581618 41826 581854
rect 42062 581618 42146 581854
rect 42382 581618 42414 581854
rect 41794 581534 42414 581618
rect 41794 581298 41826 581534
rect 42062 581298 42146 581534
rect 42382 581298 42414 581534
rect 77794 581618 77826 581854
rect 78062 581618 78146 581854
rect 78382 581618 78414 581854
rect 77794 581534 78414 581618
rect 77794 581298 77826 581534
rect 78062 581298 78146 581534
rect 78382 581298 78414 581534
rect 113794 581618 113826 581854
rect 114062 581618 114146 581854
rect 114382 581618 114414 581854
rect 113794 581534 114414 581618
rect 113794 581298 113826 581534
rect 114062 581298 114146 581534
rect 114382 581298 114414 581534
rect 149794 581618 149826 581854
rect 150062 581618 150146 581854
rect 150382 581618 150414 581854
rect 149794 581534 150414 581618
rect 149794 581298 149826 581534
rect 150062 581298 150146 581534
rect 150382 581298 150414 581534
rect 185794 581618 185826 581854
rect 186062 581618 186146 581854
rect 186382 581618 186414 581854
rect 185794 581534 186414 581618
rect 185794 581298 185826 581534
rect 186062 581298 186146 581534
rect 186382 581298 186414 581534
rect 221794 581618 221826 581854
rect 222062 581618 222146 581854
rect 222382 581618 222414 581854
rect 221794 581534 222414 581618
rect 221794 581298 221826 581534
rect 222062 581298 222146 581534
rect 222382 581298 222414 581534
rect 257794 581618 257826 581854
rect 258062 581618 258146 581854
rect 258382 581618 258414 581854
rect 257794 581534 258414 581618
rect 257794 581298 257826 581534
rect 258062 581298 258146 581534
rect 258382 581298 258414 581534
rect 293794 581618 293826 581854
rect 294062 581618 294146 581854
rect 294382 581618 294414 581854
rect 293794 581534 294414 581618
rect 293794 581298 293826 581534
rect 294062 581298 294146 581534
rect 294382 581298 294414 581534
rect 329794 581618 329826 581854
rect 330062 581618 330146 581854
rect 330382 581618 330414 581854
rect 329794 581534 330414 581618
rect 329794 581298 329826 581534
rect 330062 581298 330146 581534
rect 330382 581298 330414 581534
rect 365794 581618 365826 581854
rect 366062 581618 366146 581854
rect 366382 581618 366414 581854
rect 365794 581534 366414 581618
rect 365794 581298 365826 581534
rect 366062 581298 366146 581534
rect 366382 581298 366414 581534
rect 401794 581618 401826 581854
rect 402062 581618 402146 581854
rect 402382 581618 402414 581854
rect 401794 581534 402414 581618
rect 401794 581298 401826 581534
rect 402062 581298 402146 581534
rect 402382 581298 402414 581534
rect 437794 581618 437826 581854
rect 438062 581618 438146 581854
rect 438382 581618 438414 581854
rect 437794 581534 438414 581618
rect 437794 581298 437826 581534
rect 438062 581298 438146 581534
rect 438382 581298 438414 581534
rect 473794 581618 473826 581854
rect 474062 581618 474146 581854
rect 474382 581618 474414 581854
rect 473794 581534 474414 581618
rect 473794 581298 473826 581534
rect 474062 581298 474146 581534
rect 474382 581298 474414 581534
rect 509794 581618 509826 581854
rect 510062 581618 510146 581854
rect 510382 581618 510414 581854
rect 509794 581534 510414 581618
rect 509794 581298 509826 581534
rect 510062 581298 510146 581534
rect 510382 581298 510414 581534
rect 545794 581618 545826 581854
rect 546062 581618 546146 581854
rect 546382 581618 546414 581854
rect 545794 581534 546414 581618
rect 545794 581298 545826 581534
rect 546062 581298 546146 581534
rect 546382 581298 546414 581534
rect -2006 545854 -1386 581298
rect 582294 550354 582914 585798
rect 13166 550118 13198 550354
rect 13434 550118 13518 550354
rect 13754 550118 13786 550354
rect 13166 550034 13786 550118
rect 13166 549798 13198 550034
rect 13434 549798 13518 550034
rect 13754 549798 13786 550034
rect 167794 550118 167826 550354
rect 168062 550118 168146 550354
rect 168382 550118 168414 550354
rect 167794 550034 168414 550118
rect 167794 549798 167826 550034
rect 168062 549798 168146 550034
rect 168382 549798 168414 550034
rect 203794 550118 203826 550354
rect 204062 550118 204146 550354
rect 204382 550118 204414 550354
rect 203794 550034 204414 550118
rect 203794 549798 203826 550034
rect 204062 549798 204146 550034
rect 204382 549798 204414 550034
rect 239794 550118 239826 550354
rect 240062 550118 240146 550354
rect 240382 550118 240414 550354
rect 239794 550034 240414 550118
rect 239794 549798 239826 550034
rect 240062 549798 240146 550034
rect 240382 549798 240414 550034
rect 275794 550118 275826 550354
rect 276062 550118 276146 550354
rect 276382 550118 276414 550354
rect 275794 550034 276414 550118
rect 275794 549798 275826 550034
rect 276062 549798 276146 550034
rect 276382 549798 276414 550034
rect 311794 550118 311826 550354
rect 312062 550118 312146 550354
rect 312382 550118 312414 550354
rect 311794 550034 312414 550118
rect 311794 549798 311826 550034
rect 312062 549798 312146 550034
rect 312382 549798 312414 550034
rect 347794 550118 347826 550354
rect 348062 550118 348146 550354
rect 348382 550118 348414 550354
rect 347794 550034 348414 550118
rect 347794 549798 347826 550034
rect 348062 549798 348146 550034
rect 348382 549798 348414 550034
rect 383794 550118 383826 550354
rect 384062 550118 384146 550354
rect 384382 550118 384414 550354
rect 383794 550034 384414 550118
rect 383794 549798 383826 550034
rect 384062 549798 384146 550034
rect 384382 549798 384414 550034
rect 419794 550118 419826 550354
rect 420062 550118 420146 550354
rect 420382 550118 420414 550354
rect 419794 550034 420414 550118
rect 419794 549798 419826 550034
rect 420062 549798 420146 550034
rect 420382 549798 420414 550034
rect 563794 550118 563826 550354
rect 564062 550118 564146 550354
rect 564382 550118 564414 550354
rect 563794 550034 564414 550118
rect 563794 549798 563826 550034
rect 564062 549798 564146 550034
rect 564382 549798 564414 550034
rect 582294 550118 582326 550354
rect 582562 550118 582646 550354
rect 582882 550118 582914 550354
rect 582294 550034 582914 550118
rect 582294 549798 582326 550034
rect 582562 549798 582646 550034
rect 582882 549798 582914 550034
rect -2006 545618 -1974 545854
rect -1738 545618 -1654 545854
rect -1418 545618 -1386 545854
rect -2006 545534 -1386 545618
rect -2006 545298 -1974 545534
rect -1738 545298 -1654 545534
rect -1418 545298 -1386 545534
rect 5794 545618 5826 545854
rect 6062 545618 6146 545854
rect 6382 545618 6414 545854
rect 5794 545534 6414 545618
rect 5794 545298 5826 545534
rect 6062 545298 6146 545534
rect 6382 545298 6414 545534
rect 185794 545618 185826 545854
rect 186062 545618 186146 545854
rect 186382 545618 186414 545854
rect 185794 545534 186414 545618
rect 185794 545298 185826 545534
rect 186062 545298 186146 545534
rect 186382 545298 186414 545534
rect 221794 545618 221826 545854
rect 222062 545618 222146 545854
rect 222382 545618 222414 545854
rect 221794 545534 222414 545618
rect 221794 545298 221826 545534
rect 222062 545298 222146 545534
rect 222382 545298 222414 545534
rect 257794 545618 257826 545854
rect 258062 545618 258146 545854
rect 258382 545618 258414 545854
rect 257794 545534 258414 545618
rect 257794 545298 257826 545534
rect 258062 545298 258146 545534
rect 258382 545298 258414 545534
rect 293794 545618 293826 545854
rect 294062 545618 294146 545854
rect 294382 545618 294414 545854
rect 293794 545534 294414 545618
rect 293794 545298 293826 545534
rect 294062 545298 294146 545534
rect 294382 545298 294414 545534
rect 329794 545618 329826 545854
rect 330062 545618 330146 545854
rect 330382 545618 330414 545854
rect 329794 545534 330414 545618
rect 329794 545298 329826 545534
rect 330062 545298 330146 545534
rect 330382 545298 330414 545534
rect 365794 545618 365826 545854
rect 366062 545618 366146 545854
rect 366382 545618 366414 545854
rect 365794 545534 366414 545618
rect 365794 545298 365826 545534
rect 366062 545298 366146 545534
rect 366382 545298 366414 545534
rect 401794 545618 401826 545854
rect 402062 545618 402146 545854
rect 402382 545618 402414 545854
rect 401794 545534 402414 545618
rect 401794 545298 401826 545534
rect 402062 545298 402146 545534
rect 402382 545298 402414 545534
rect 570318 545618 570350 545854
rect 570586 545618 570670 545854
rect 570906 545618 570938 545854
rect 570318 545534 570938 545618
rect 570318 545298 570350 545534
rect 570586 545298 570670 545534
rect 570906 545298 570938 545534
rect -2006 509854 -1386 545298
rect 582294 514354 582914 549798
rect 13166 514118 13198 514354
rect 13434 514118 13518 514354
rect 13754 514118 13786 514354
rect 13166 514034 13786 514118
rect 13166 513798 13198 514034
rect 13434 513798 13518 514034
rect 13754 513798 13786 514034
rect 167794 514118 167826 514354
rect 168062 514118 168146 514354
rect 168382 514118 168414 514354
rect 167794 514034 168414 514118
rect 167794 513798 167826 514034
rect 168062 513798 168146 514034
rect 168382 513798 168414 514034
rect 203794 514118 203826 514354
rect 204062 514118 204146 514354
rect 204382 514118 204414 514354
rect 203794 514034 204414 514118
rect 203794 513798 203826 514034
rect 204062 513798 204146 514034
rect 204382 513798 204414 514034
rect 239794 514118 239826 514354
rect 240062 514118 240146 514354
rect 240382 514118 240414 514354
rect 239794 514034 240414 514118
rect 239794 513798 239826 514034
rect 240062 513798 240146 514034
rect 240382 513798 240414 514034
rect 275794 514118 275826 514354
rect 276062 514118 276146 514354
rect 276382 514118 276414 514354
rect 275794 514034 276414 514118
rect 275794 513798 275826 514034
rect 276062 513798 276146 514034
rect 276382 513798 276414 514034
rect 311794 514118 311826 514354
rect 312062 514118 312146 514354
rect 312382 514118 312414 514354
rect 311794 514034 312414 514118
rect 311794 513798 311826 514034
rect 312062 513798 312146 514034
rect 312382 513798 312414 514034
rect 347794 514118 347826 514354
rect 348062 514118 348146 514354
rect 348382 514118 348414 514354
rect 347794 514034 348414 514118
rect 347794 513798 347826 514034
rect 348062 513798 348146 514034
rect 348382 513798 348414 514034
rect 383794 514118 383826 514354
rect 384062 514118 384146 514354
rect 384382 514118 384414 514354
rect 383794 514034 384414 514118
rect 383794 513798 383826 514034
rect 384062 513798 384146 514034
rect 384382 513798 384414 514034
rect 419794 514118 419826 514354
rect 420062 514118 420146 514354
rect 420382 514118 420414 514354
rect 419794 514034 420414 514118
rect 419794 513798 419826 514034
rect 420062 513798 420146 514034
rect 420382 513798 420414 514034
rect 563794 514118 563826 514354
rect 564062 514118 564146 514354
rect 564382 514118 564414 514354
rect 563794 514034 564414 514118
rect 563794 513798 563826 514034
rect 564062 513798 564146 514034
rect 564382 513798 564414 514034
rect 582294 514118 582326 514354
rect 582562 514118 582646 514354
rect 582882 514118 582914 514354
rect 582294 514034 582914 514118
rect 582294 513798 582326 514034
rect 582562 513798 582646 514034
rect 582882 513798 582914 514034
rect -2006 509618 -1974 509854
rect -1738 509618 -1654 509854
rect -1418 509618 -1386 509854
rect -2006 509534 -1386 509618
rect -2006 509298 -1974 509534
rect -1738 509298 -1654 509534
rect -1418 509298 -1386 509534
rect 5794 509618 5826 509854
rect 6062 509618 6146 509854
rect 6382 509618 6414 509854
rect 5794 509534 6414 509618
rect 5794 509298 5826 509534
rect 6062 509298 6146 509534
rect 6382 509298 6414 509534
rect 185794 509618 185826 509854
rect 186062 509618 186146 509854
rect 186382 509618 186414 509854
rect 185794 509534 186414 509618
rect 185794 509298 185826 509534
rect 186062 509298 186146 509534
rect 186382 509298 186414 509534
rect 221794 509618 221826 509854
rect 222062 509618 222146 509854
rect 222382 509618 222414 509854
rect 221794 509534 222414 509618
rect 221794 509298 221826 509534
rect 222062 509298 222146 509534
rect 222382 509298 222414 509534
rect 257794 509618 257826 509854
rect 258062 509618 258146 509854
rect 258382 509618 258414 509854
rect 257794 509534 258414 509618
rect 257794 509298 257826 509534
rect 258062 509298 258146 509534
rect 258382 509298 258414 509534
rect 293794 509618 293826 509854
rect 294062 509618 294146 509854
rect 294382 509618 294414 509854
rect 293794 509534 294414 509618
rect 293794 509298 293826 509534
rect 294062 509298 294146 509534
rect 294382 509298 294414 509534
rect 329794 509618 329826 509854
rect 330062 509618 330146 509854
rect 330382 509618 330414 509854
rect 329794 509534 330414 509618
rect 329794 509298 329826 509534
rect 330062 509298 330146 509534
rect 330382 509298 330414 509534
rect 365794 509618 365826 509854
rect 366062 509618 366146 509854
rect 366382 509618 366414 509854
rect 365794 509534 366414 509618
rect 365794 509298 365826 509534
rect 366062 509298 366146 509534
rect 366382 509298 366414 509534
rect 401794 509618 401826 509854
rect 402062 509618 402146 509854
rect 402382 509618 402414 509854
rect 401794 509534 402414 509618
rect 401794 509298 401826 509534
rect 402062 509298 402146 509534
rect 402382 509298 402414 509534
rect 570318 509618 570350 509854
rect 570586 509618 570670 509854
rect 570906 509618 570938 509854
rect 570318 509534 570938 509618
rect 570318 509298 570350 509534
rect 570586 509298 570670 509534
rect 570906 509298 570938 509534
rect -2006 473854 -1386 509298
rect 582294 478354 582914 513798
rect 23794 478118 23826 478354
rect 24062 478118 24146 478354
rect 24382 478118 24414 478354
rect 23794 478034 24414 478118
rect 23794 477798 23826 478034
rect 24062 477798 24146 478034
rect 24382 477798 24414 478034
rect 59794 478118 59826 478354
rect 60062 478118 60146 478354
rect 60382 478118 60414 478354
rect 59794 478034 60414 478118
rect 59794 477798 59826 478034
rect 60062 477798 60146 478034
rect 60382 477798 60414 478034
rect 95794 478118 95826 478354
rect 96062 478118 96146 478354
rect 96382 478118 96414 478354
rect 95794 478034 96414 478118
rect 95794 477798 95826 478034
rect 96062 477798 96146 478034
rect 96382 477798 96414 478034
rect 131794 478118 131826 478354
rect 132062 478118 132146 478354
rect 132382 478118 132414 478354
rect 131794 478034 132414 478118
rect 131794 477798 131826 478034
rect 132062 477798 132146 478034
rect 132382 477798 132414 478034
rect 167794 478118 167826 478354
rect 168062 478118 168146 478354
rect 168382 478118 168414 478354
rect 167794 478034 168414 478118
rect 167794 477798 167826 478034
rect 168062 477798 168146 478034
rect 168382 477798 168414 478034
rect 203794 478118 203826 478354
rect 204062 478118 204146 478354
rect 204382 478118 204414 478354
rect 203794 478034 204414 478118
rect 203794 477798 203826 478034
rect 204062 477798 204146 478034
rect 204382 477798 204414 478034
rect 239794 478118 239826 478354
rect 240062 478118 240146 478354
rect 240382 478118 240414 478354
rect 239794 478034 240414 478118
rect 239794 477798 239826 478034
rect 240062 477798 240146 478034
rect 240382 477798 240414 478034
rect 275794 478118 275826 478354
rect 276062 478118 276146 478354
rect 276382 478118 276414 478354
rect 275794 478034 276414 478118
rect 275794 477798 275826 478034
rect 276062 477798 276146 478034
rect 276382 477798 276414 478034
rect 311794 478118 311826 478354
rect 312062 478118 312146 478354
rect 312382 478118 312414 478354
rect 311794 478034 312414 478118
rect 311794 477798 311826 478034
rect 312062 477798 312146 478034
rect 312382 477798 312414 478034
rect 347794 478118 347826 478354
rect 348062 478118 348146 478354
rect 348382 478118 348414 478354
rect 347794 478034 348414 478118
rect 347794 477798 347826 478034
rect 348062 477798 348146 478034
rect 348382 477798 348414 478034
rect 383794 478118 383826 478354
rect 384062 478118 384146 478354
rect 384382 478118 384414 478354
rect 383794 478034 384414 478118
rect 383794 477798 383826 478034
rect 384062 477798 384146 478034
rect 384382 477798 384414 478034
rect 419794 478118 419826 478354
rect 420062 478118 420146 478354
rect 420382 478118 420414 478354
rect 419794 478034 420414 478118
rect 419794 477798 419826 478034
rect 420062 477798 420146 478034
rect 420382 477798 420414 478034
rect 455794 478118 455826 478354
rect 456062 478118 456146 478354
rect 456382 478118 456414 478354
rect 455794 478034 456414 478118
rect 455794 477798 455826 478034
rect 456062 477798 456146 478034
rect 456382 477798 456414 478034
rect 491794 478118 491826 478354
rect 492062 478118 492146 478354
rect 492382 478118 492414 478354
rect 491794 478034 492414 478118
rect 491794 477798 491826 478034
rect 492062 477798 492146 478034
rect 492382 477798 492414 478034
rect 527794 478118 527826 478354
rect 528062 478118 528146 478354
rect 528382 478118 528414 478354
rect 527794 478034 528414 478118
rect 527794 477798 527826 478034
rect 528062 477798 528146 478034
rect 528382 477798 528414 478034
rect 563794 478118 563826 478354
rect 564062 478118 564146 478354
rect 564382 478118 564414 478354
rect 563794 478034 564414 478118
rect 563794 477798 563826 478034
rect 564062 477798 564146 478034
rect 564382 477798 564414 478034
rect 582294 478118 582326 478354
rect 582562 478118 582646 478354
rect 582882 478118 582914 478354
rect 582294 478034 582914 478118
rect 582294 477798 582326 478034
rect 582562 477798 582646 478034
rect 582882 477798 582914 478034
rect -2006 473618 -1974 473854
rect -1738 473618 -1654 473854
rect -1418 473618 -1386 473854
rect -2006 473534 -1386 473618
rect -2006 473298 -1974 473534
rect -1738 473298 -1654 473534
rect -1418 473298 -1386 473534
rect 5794 473618 5826 473854
rect 6062 473618 6146 473854
rect 6382 473618 6414 473854
rect 5794 473534 6414 473618
rect 5794 473298 5826 473534
rect 6062 473298 6146 473534
rect 6382 473298 6414 473534
rect 41794 473618 41826 473854
rect 42062 473618 42146 473854
rect 42382 473618 42414 473854
rect 41794 473534 42414 473618
rect 41794 473298 41826 473534
rect 42062 473298 42146 473534
rect 42382 473298 42414 473534
rect 77794 473618 77826 473854
rect 78062 473618 78146 473854
rect 78382 473618 78414 473854
rect 77794 473534 78414 473618
rect 77794 473298 77826 473534
rect 78062 473298 78146 473534
rect 78382 473298 78414 473534
rect 113794 473618 113826 473854
rect 114062 473618 114146 473854
rect 114382 473618 114414 473854
rect 113794 473534 114414 473618
rect 113794 473298 113826 473534
rect 114062 473298 114146 473534
rect 114382 473298 114414 473534
rect 149794 473618 149826 473854
rect 150062 473618 150146 473854
rect 150382 473618 150414 473854
rect 149794 473534 150414 473618
rect 149794 473298 149826 473534
rect 150062 473298 150146 473534
rect 150382 473298 150414 473534
rect 185794 473618 185826 473854
rect 186062 473618 186146 473854
rect 186382 473618 186414 473854
rect 185794 473534 186414 473618
rect 185794 473298 185826 473534
rect 186062 473298 186146 473534
rect 186382 473298 186414 473534
rect 221794 473618 221826 473854
rect 222062 473618 222146 473854
rect 222382 473618 222414 473854
rect 221794 473534 222414 473618
rect 221794 473298 221826 473534
rect 222062 473298 222146 473534
rect 222382 473298 222414 473534
rect 257794 473618 257826 473854
rect 258062 473618 258146 473854
rect 258382 473618 258414 473854
rect 257794 473534 258414 473618
rect 257794 473298 257826 473534
rect 258062 473298 258146 473534
rect 258382 473298 258414 473534
rect 293794 473618 293826 473854
rect 294062 473618 294146 473854
rect 294382 473618 294414 473854
rect 293794 473534 294414 473618
rect 293794 473298 293826 473534
rect 294062 473298 294146 473534
rect 294382 473298 294414 473534
rect 329794 473618 329826 473854
rect 330062 473618 330146 473854
rect 330382 473618 330414 473854
rect 329794 473534 330414 473618
rect 329794 473298 329826 473534
rect 330062 473298 330146 473534
rect 330382 473298 330414 473534
rect 365794 473618 365826 473854
rect 366062 473618 366146 473854
rect 366382 473618 366414 473854
rect 365794 473534 366414 473618
rect 365794 473298 365826 473534
rect 366062 473298 366146 473534
rect 366382 473298 366414 473534
rect 401794 473618 401826 473854
rect 402062 473618 402146 473854
rect 402382 473618 402414 473854
rect 401794 473534 402414 473618
rect 401794 473298 401826 473534
rect 402062 473298 402146 473534
rect 402382 473298 402414 473534
rect 437794 473618 437826 473854
rect 438062 473618 438146 473854
rect 438382 473618 438414 473854
rect 437794 473534 438414 473618
rect 437794 473298 437826 473534
rect 438062 473298 438146 473534
rect 438382 473298 438414 473534
rect 473794 473618 473826 473854
rect 474062 473618 474146 473854
rect 474382 473618 474414 473854
rect 473794 473534 474414 473618
rect 473794 473298 473826 473534
rect 474062 473298 474146 473534
rect 474382 473298 474414 473534
rect 509794 473618 509826 473854
rect 510062 473618 510146 473854
rect 510382 473618 510414 473854
rect 509794 473534 510414 473618
rect 509794 473298 509826 473534
rect 510062 473298 510146 473534
rect 510382 473298 510414 473534
rect 545794 473618 545826 473854
rect 546062 473618 546146 473854
rect 546382 473618 546414 473854
rect 545794 473534 546414 473618
rect 545794 473298 545826 473534
rect 546062 473298 546146 473534
rect 546382 473298 546414 473534
rect -2006 437854 -1386 473298
rect 582294 442354 582914 477798
rect 13166 442118 13198 442354
rect 13434 442118 13518 442354
rect 13754 442118 13786 442354
rect 13166 442034 13786 442118
rect 13166 441798 13198 442034
rect 13434 441798 13518 442034
rect 13754 441798 13786 442034
rect 167794 442118 167826 442354
rect 168062 442118 168146 442354
rect 168382 442118 168414 442354
rect 167794 442034 168414 442118
rect 167794 441798 167826 442034
rect 168062 441798 168146 442034
rect 168382 441798 168414 442034
rect 203794 442118 203826 442354
rect 204062 442118 204146 442354
rect 204382 442118 204414 442354
rect 203794 442034 204414 442118
rect 203794 441798 203826 442034
rect 204062 441798 204146 442034
rect 204382 441798 204414 442034
rect 239794 442118 239826 442354
rect 240062 442118 240146 442354
rect 240382 442118 240414 442354
rect 239794 442034 240414 442118
rect 239794 441798 239826 442034
rect 240062 441798 240146 442034
rect 240382 441798 240414 442034
rect 275794 442118 275826 442354
rect 276062 442118 276146 442354
rect 276382 442118 276414 442354
rect 275794 442034 276414 442118
rect 275794 441798 275826 442034
rect 276062 441798 276146 442034
rect 276382 441798 276414 442034
rect 311794 442118 311826 442354
rect 312062 442118 312146 442354
rect 312382 442118 312414 442354
rect 311794 442034 312414 442118
rect 311794 441798 311826 442034
rect 312062 441798 312146 442034
rect 312382 441798 312414 442034
rect 347794 442118 347826 442354
rect 348062 442118 348146 442354
rect 348382 442118 348414 442354
rect 347794 442034 348414 442118
rect 347794 441798 347826 442034
rect 348062 441798 348146 442034
rect 348382 441798 348414 442034
rect 383794 442118 383826 442354
rect 384062 442118 384146 442354
rect 384382 442118 384414 442354
rect 383794 442034 384414 442118
rect 383794 441798 383826 442034
rect 384062 441798 384146 442034
rect 384382 441798 384414 442034
rect 419794 442118 419826 442354
rect 420062 442118 420146 442354
rect 420382 442118 420414 442354
rect 419794 442034 420414 442118
rect 419794 441798 419826 442034
rect 420062 441798 420146 442034
rect 420382 441798 420414 442034
rect 563794 442118 563826 442354
rect 564062 442118 564146 442354
rect 564382 442118 564414 442354
rect 563794 442034 564414 442118
rect 563794 441798 563826 442034
rect 564062 441798 564146 442034
rect 564382 441798 564414 442034
rect 582294 442118 582326 442354
rect 582562 442118 582646 442354
rect 582882 442118 582914 442354
rect 582294 442034 582914 442118
rect 582294 441798 582326 442034
rect 582562 441798 582646 442034
rect 582882 441798 582914 442034
rect -2006 437618 -1974 437854
rect -1738 437618 -1654 437854
rect -1418 437618 -1386 437854
rect -2006 437534 -1386 437618
rect -2006 437298 -1974 437534
rect -1738 437298 -1654 437534
rect -1418 437298 -1386 437534
rect 5794 437618 5826 437854
rect 6062 437618 6146 437854
rect 6382 437618 6414 437854
rect 5794 437534 6414 437618
rect 5794 437298 5826 437534
rect 6062 437298 6146 437534
rect 6382 437298 6414 437534
rect 185794 437618 185826 437854
rect 186062 437618 186146 437854
rect 186382 437618 186414 437854
rect 185794 437534 186414 437618
rect 185794 437298 185826 437534
rect 186062 437298 186146 437534
rect 186382 437298 186414 437534
rect 221794 437618 221826 437854
rect 222062 437618 222146 437854
rect 222382 437618 222414 437854
rect 221794 437534 222414 437618
rect 221794 437298 221826 437534
rect 222062 437298 222146 437534
rect 222382 437298 222414 437534
rect 257794 437618 257826 437854
rect 258062 437618 258146 437854
rect 258382 437618 258414 437854
rect 257794 437534 258414 437618
rect 257794 437298 257826 437534
rect 258062 437298 258146 437534
rect 258382 437298 258414 437534
rect 293794 437618 293826 437854
rect 294062 437618 294146 437854
rect 294382 437618 294414 437854
rect 293794 437534 294414 437618
rect 293794 437298 293826 437534
rect 294062 437298 294146 437534
rect 294382 437298 294414 437534
rect 329794 437618 329826 437854
rect 330062 437618 330146 437854
rect 330382 437618 330414 437854
rect 329794 437534 330414 437618
rect 329794 437298 329826 437534
rect 330062 437298 330146 437534
rect 330382 437298 330414 437534
rect 365794 437618 365826 437854
rect 366062 437618 366146 437854
rect 366382 437618 366414 437854
rect 365794 437534 366414 437618
rect 365794 437298 365826 437534
rect 366062 437298 366146 437534
rect 366382 437298 366414 437534
rect 401794 437618 401826 437854
rect 402062 437618 402146 437854
rect 402382 437618 402414 437854
rect 401794 437534 402414 437618
rect 401794 437298 401826 437534
rect 402062 437298 402146 437534
rect 402382 437298 402414 437534
rect 570318 437618 570350 437854
rect 570586 437618 570670 437854
rect 570906 437618 570938 437854
rect 570318 437534 570938 437618
rect 570318 437298 570350 437534
rect 570586 437298 570670 437534
rect 570906 437298 570938 437534
rect -2006 401854 -1386 437298
rect 582294 406354 582914 441798
rect 13166 406118 13198 406354
rect 13434 406118 13518 406354
rect 13754 406118 13786 406354
rect 13166 406034 13786 406118
rect 13166 405798 13198 406034
rect 13434 405798 13518 406034
rect 13754 405798 13786 406034
rect 167794 406118 167826 406354
rect 168062 406118 168146 406354
rect 168382 406118 168414 406354
rect 167794 406034 168414 406118
rect 167794 405798 167826 406034
rect 168062 405798 168146 406034
rect 168382 405798 168414 406034
rect 203794 406118 203826 406354
rect 204062 406118 204146 406354
rect 204382 406118 204414 406354
rect 203794 406034 204414 406118
rect 203794 405798 203826 406034
rect 204062 405798 204146 406034
rect 204382 405798 204414 406034
rect 239794 406118 239826 406354
rect 240062 406118 240146 406354
rect 240382 406118 240414 406354
rect 239794 406034 240414 406118
rect 239794 405798 239826 406034
rect 240062 405798 240146 406034
rect 240382 405798 240414 406034
rect 275794 406118 275826 406354
rect 276062 406118 276146 406354
rect 276382 406118 276414 406354
rect 275794 406034 276414 406118
rect 275794 405798 275826 406034
rect 276062 405798 276146 406034
rect 276382 405798 276414 406034
rect 311794 406118 311826 406354
rect 312062 406118 312146 406354
rect 312382 406118 312414 406354
rect 311794 406034 312414 406118
rect 311794 405798 311826 406034
rect 312062 405798 312146 406034
rect 312382 405798 312414 406034
rect 347794 406118 347826 406354
rect 348062 406118 348146 406354
rect 348382 406118 348414 406354
rect 347794 406034 348414 406118
rect 347794 405798 347826 406034
rect 348062 405798 348146 406034
rect 348382 405798 348414 406034
rect 383794 406118 383826 406354
rect 384062 406118 384146 406354
rect 384382 406118 384414 406354
rect 383794 406034 384414 406118
rect 383794 405798 383826 406034
rect 384062 405798 384146 406034
rect 384382 405798 384414 406034
rect 419794 406118 419826 406354
rect 420062 406118 420146 406354
rect 420382 406118 420414 406354
rect 419794 406034 420414 406118
rect 419794 405798 419826 406034
rect 420062 405798 420146 406034
rect 420382 405798 420414 406034
rect 563794 406118 563826 406354
rect 564062 406118 564146 406354
rect 564382 406118 564414 406354
rect 563794 406034 564414 406118
rect 563794 405798 563826 406034
rect 564062 405798 564146 406034
rect 564382 405798 564414 406034
rect 582294 406118 582326 406354
rect 582562 406118 582646 406354
rect 582882 406118 582914 406354
rect 582294 406034 582914 406118
rect 582294 405798 582326 406034
rect 582562 405798 582646 406034
rect 582882 405798 582914 406034
rect -2006 401618 -1974 401854
rect -1738 401618 -1654 401854
rect -1418 401618 -1386 401854
rect -2006 401534 -1386 401618
rect -2006 401298 -1974 401534
rect -1738 401298 -1654 401534
rect -1418 401298 -1386 401534
rect 5794 401618 5826 401854
rect 6062 401618 6146 401854
rect 6382 401618 6414 401854
rect 5794 401534 6414 401618
rect 5794 401298 5826 401534
rect 6062 401298 6146 401534
rect 6382 401298 6414 401534
rect 185794 401618 185826 401854
rect 186062 401618 186146 401854
rect 186382 401618 186414 401854
rect 185794 401534 186414 401618
rect 185794 401298 185826 401534
rect 186062 401298 186146 401534
rect 186382 401298 186414 401534
rect 221794 401618 221826 401854
rect 222062 401618 222146 401854
rect 222382 401618 222414 401854
rect 221794 401534 222414 401618
rect 221794 401298 221826 401534
rect 222062 401298 222146 401534
rect 222382 401298 222414 401534
rect 257794 401618 257826 401854
rect 258062 401618 258146 401854
rect 258382 401618 258414 401854
rect 257794 401534 258414 401618
rect 257794 401298 257826 401534
rect 258062 401298 258146 401534
rect 258382 401298 258414 401534
rect 293794 401618 293826 401854
rect 294062 401618 294146 401854
rect 294382 401618 294414 401854
rect 293794 401534 294414 401618
rect 293794 401298 293826 401534
rect 294062 401298 294146 401534
rect 294382 401298 294414 401534
rect 329794 401618 329826 401854
rect 330062 401618 330146 401854
rect 330382 401618 330414 401854
rect 329794 401534 330414 401618
rect 329794 401298 329826 401534
rect 330062 401298 330146 401534
rect 330382 401298 330414 401534
rect 365794 401618 365826 401854
rect 366062 401618 366146 401854
rect 366382 401618 366414 401854
rect 365794 401534 366414 401618
rect 365794 401298 365826 401534
rect 366062 401298 366146 401534
rect 366382 401298 366414 401534
rect 401794 401618 401826 401854
rect 402062 401618 402146 401854
rect 402382 401618 402414 401854
rect 401794 401534 402414 401618
rect 401794 401298 401826 401534
rect 402062 401298 402146 401534
rect 402382 401298 402414 401534
rect 570318 401618 570350 401854
rect 570586 401618 570670 401854
rect 570906 401618 570938 401854
rect 570318 401534 570938 401618
rect 570318 401298 570350 401534
rect 570586 401298 570670 401534
rect 570906 401298 570938 401534
rect -2006 365854 -1386 401298
rect 582294 370354 582914 405798
rect 13166 370118 13198 370354
rect 13434 370118 13518 370354
rect 13754 370118 13786 370354
rect 13166 370034 13786 370118
rect 13166 369798 13198 370034
rect 13434 369798 13518 370034
rect 13754 369798 13786 370034
rect 167794 370118 167826 370354
rect 168062 370118 168146 370354
rect 168382 370118 168414 370354
rect 167794 370034 168414 370118
rect 167794 369798 167826 370034
rect 168062 369798 168146 370034
rect 168382 369798 168414 370034
rect 203794 370118 203826 370354
rect 204062 370118 204146 370354
rect 204382 370118 204414 370354
rect 203794 370034 204414 370118
rect 203794 369798 203826 370034
rect 204062 369798 204146 370034
rect 204382 369798 204414 370034
rect 239794 370118 239826 370354
rect 240062 370118 240146 370354
rect 240382 370118 240414 370354
rect 239794 370034 240414 370118
rect 239794 369798 239826 370034
rect 240062 369798 240146 370034
rect 240382 369798 240414 370034
rect 275794 370118 275826 370354
rect 276062 370118 276146 370354
rect 276382 370118 276414 370354
rect 275794 370034 276414 370118
rect 275794 369798 275826 370034
rect 276062 369798 276146 370034
rect 276382 369798 276414 370034
rect 311794 370118 311826 370354
rect 312062 370118 312146 370354
rect 312382 370118 312414 370354
rect 311794 370034 312414 370118
rect 311794 369798 311826 370034
rect 312062 369798 312146 370034
rect 312382 369798 312414 370034
rect 347794 370118 347826 370354
rect 348062 370118 348146 370354
rect 348382 370118 348414 370354
rect 347794 370034 348414 370118
rect 347794 369798 347826 370034
rect 348062 369798 348146 370034
rect 348382 369798 348414 370034
rect 383794 370118 383826 370354
rect 384062 370118 384146 370354
rect 384382 370118 384414 370354
rect 383794 370034 384414 370118
rect 383794 369798 383826 370034
rect 384062 369798 384146 370034
rect 384382 369798 384414 370034
rect 419794 370118 419826 370354
rect 420062 370118 420146 370354
rect 420382 370118 420414 370354
rect 419794 370034 420414 370118
rect 419794 369798 419826 370034
rect 420062 369798 420146 370034
rect 420382 369798 420414 370034
rect 563794 370118 563826 370354
rect 564062 370118 564146 370354
rect 564382 370118 564414 370354
rect 563794 370034 564414 370118
rect 563794 369798 563826 370034
rect 564062 369798 564146 370034
rect 564382 369798 564414 370034
rect 582294 370118 582326 370354
rect 582562 370118 582646 370354
rect 582882 370118 582914 370354
rect 582294 370034 582914 370118
rect 582294 369798 582326 370034
rect 582562 369798 582646 370034
rect 582882 369798 582914 370034
rect -2006 365618 -1974 365854
rect -1738 365618 -1654 365854
rect -1418 365618 -1386 365854
rect -2006 365534 -1386 365618
rect -2006 365298 -1974 365534
rect -1738 365298 -1654 365534
rect -1418 365298 -1386 365534
rect 5794 365618 5826 365854
rect 6062 365618 6146 365854
rect 6382 365618 6414 365854
rect 5794 365534 6414 365618
rect 5794 365298 5826 365534
rect 6062 365298 6146 365534
rect 6382 365298 6414 365534
rect 41794 365618 41826 365854
rect 42062 365618 42146 365854
rect 42382 365618 42414 365854
rect 41794 365534 42414 365618
rect 41794 365298 41826 365534
rect 42062 365298 42146 365534
rect 42382 365298 42414 365534
rect 77794 365618 77826 365854
rect 78062 365618 78146 365854
rect 78382 365618 78414 365854
rect 77794 365534 78414 365618
rect 77794 365298 77826 365534
rect 78062 365298 78146 365534
rect 78382 365298 78414 365534
rect 113794 365618 113826 365854
rect 114062 365618 114146 365854
rect 114382 365618 114414 365854
rect 113794 365534 114414 365618
rect 113794 365298 113826 365534
rect 114062 365298 114146 365534
rect 114382 365298 114414 365534
rect 149794 365618 149826 365854
rect 150062 365618 150146 365854
rect 150382 365618 150414 365854
rect 149794 365534 150414 365618
rect 149794 365298 149826 365534
rect 150062 365298 150146 365534
rect 150382 365298 150414 365534
rect 185794 365618 185826 365854
rect 186062 365618 186146 365854
rect 186382 365618 186414 365854
rect 185794 365534 186414 365618
rect 185794 365298 185826 365534
rect 186062 365298 186146 365534
rect 186382 365298 186414 365534
rect 221794 365618 221826 365854
rect 222062 365618 222146 365854
rect 222382 365618 222414 365854
rect 221794 365534 222414 365618
rect 221794 365298 221826 365534
rect 222062 365298 222146 365534
rect 222382 365298 222414 365534
rect 257794 365618 257826 365854
rect 258062 365618 258146 365854
rect 258382 365618 258414 365854
rect 257794 365534 258414 365618
rect 257794 365298 257826 365534
rect 258062 365298 258146 365534
rect 258382 365298 258414 365534
rect 293794 365618 293826 365854
rect 294062 365618 294146 365854
rect 294382 365618 294414 365854
rect 293794 365534 294414 365618
rect 293794 365298 293826 365534
rect 294062 365298 294146 365534
rect 294382 365298 294414 365534
rect 329794 365618 329826 365854
rect 330062 365618 330146 365854
rect 330382 365618 330414 365854
rect 329794 365534 330414 365618
rect 329794 365298 329826 365534
rect 330062 365298 330146 365534
rect 330382 365298 330414 365534
rect 365794 365618 365826 365854
rect 366062 365618 366146 365854
rect 366382 365618 366414 365854
rect 365794 365534 366414 365618
rect 365794 365298 365826 365534
rect 366062 365298 366146 365534
rect 366382 365298 366414 365534
rect 401794 365618 401826 365854
rect 402062 365618 402146 365854
rect 402382 365618 402414 365854
rect 401794 365534 402414 365618
rect 401794 365298 401826 365534
rect 402062 365298 402146 365534
rect 402382 365298 402414 365534
rect 437794 365618 437826 365854
rect 438062 365618 438146 365854
rect 438382 365618 438414 365854
rect 437794 365534 438414 365618
rect 437794 365298 437826 365534
rect 438062 365298 438146 365534
rect 438382 365298 438414 365534
rect 473794 365618 473826 365854
rect 474062 365618 474146 365854
rect 474382 365618 474414 365854
rect 473794 365534 474414 365618
rect 473794 365298 473826 365534
rect 474062 365298 474146 365534
rect 474382 365298 474414 365534
rect 509794 365618 509826 365854
rect 510062 365618 510146 365854
rect 510382 365618 510414 365854
rect 509794 365534 510414 365618
rect 509794 365298 509826 365534
rect 510062 365298 510146 365534
rect 510382 365298 510414 365534
rect 545794 365618 545826 365854
rect 546062 365618 546146 365854
rect 546382 365618 546414 365854
rect 545794 365534 546414 365618
rect 545794 365298 545826 365534
rect 546062 365298 546146 365534
rect 546382 365298 546414 365534
rect -2006 329854 -1386 365298
rect 582294 334354 582914 369798
rect 13166 334118 13198 334354
rect 13434 334118 13518 334354
rect 13754 334118 13786 334354
rect 13166 334034 13786 334118
rect 13166 333798 13198 334034
rect 13434 333798 13518 334034
rect 13754 333798 13786 334034
rect 167794 334118 167826 334354
rect 168062 334118 168146 334354
rect 168382 334118 168414 334354
rect 167794 334034 168414 334118
rect 167794 333798 167826 334034
rect 168062 333798 168146 334034
rect 168382 333798 168414 334034
rect 203794 334118 203826 334354
rect 204062 334118 204146 334354
rect 204382 334118 204414 334354
rect 203794 334034 204414 334118
rect 203794 333798 203826 334034
rect 204062 333798 204146 334034
rect 204382 333798 204414 334034
rect 239794 334118 239826 334354
rect 240062 334118 240146 334354
rect 240382 334118 240414 334354
rect 239794 334034 240414 334118
rect 239794 333798 239826 334034
rect 240062 333798 240146 334034
rect 240382 333798 240414 334034
rect 275794 334118 275826 334354
rect 276062 334118 276146 334354
rect 276382 334118 276414 334354
rect 275794 334034 276414 334118
rect 275794 333798 275826 334034
rect 276062 333798 276146 334034
rect 276382 333798 276414 334034
rect 311794 334118 311826 334354
rect 312062 334118 312146 334354
rect 312382 334118 312414 334354
rect 311794 334034 312414 334118
rect 311794 333798 311826 334034
rect 312062 333798 312146 334034
rect 312382 333798 312414 334034
rect 347794 334118 347826 334354
rect 348062 334118 348146 334354
rect 348382 334118 348414 334354
rect 347794 334034 348414 334118
rect 347794 333798 347826 334034
rect 348062 333798 348146 334034
rect 348382 333798 348414 334034
rect 383794 334118 383826 334354
rect 384062 334118 384146 334354
rect 384382 334118 384414 334354
rect 383794 334034 384414 334118
rect 383794 333798 383826 334034
rect 384062 333798 384146 334034
rect 384382 333798 384414 334034
rect 419794 334118 419826 334354
rect 420062 334118 420146 334354
rect 420382 334118 420414 334354
rect 419794 334034 420414 334118
rect 419794 333798 419826 334034
rect 420062 333798 420146 334034
rect 420382 333798 420414 334034
rect 563794 334118 563826 334354
rect 564062 334118 564146 334354
rect 564382 334118 564414 334354
rect 563794 334034 564414 334118
rect 563794 333798 563826 334034
rect 564062 333798 564146 334034
rect 564382 333798 564414 334034
rect 582294 334118 582326 334354
rect 582562 334118 582646 334354
rect 582882 334118 582914 334354
rect 582294 334034 582914 334118
rect 582294 333798 582326 334034
rect 582562 333798 582646 334034
rect 582882 333798 582914 334034
rect -2006 329618 -1974 329854
rect -1738 329618 -1654 329854
rect -1418 329618 -1386 329854
rect -2006 329534 -1386 329618
rect -2006 329298 -1974 329534
rect -1738 329298 -1654 329534
rect -1418 329298 -1386 329534
rect 5794 329618 5826 329854
rect 6062 329618 6146 329854
rect 6382 329618 6414 329854
rect 5794 329534 6414 329618
rect 5794 329298 5826 329534
rect 6062 329298 6146 329534
rect 6382 329298 6414 329534
rect 185794 329618 185826 329854
rect 186062 329618 186146 329854
rect 186382 329618 186414 329854
rect 185794 329534 186414 329618
rect 185794 329298 185826 329534
rect 186062 329298 186146 329534
rect 186382 329298 186414 329534
rect 221794 329618 221826 329854
rect 222062 329618 222146 329854
rect 222382 329618 222414 329854
rect 221794 329534 222414 329618
rect 221794 329298 221826 329534
rect 222062 329298 222146 329534
rect 222382 329298 222414 329534
rect 257794 329618 257826 329854
rect 258062 329618 258146 329854
rect 258382 329618 258414 329854
rect 257794 329534 258414 329618
rect 257794 329298 257826 329534
rect 258062 329298 258146 329534
rect 258382 329298 258414 329534
rect 293794 329618 293826 329854
rect 294062 329618 294146 329854
rect 294382 329618 294414 329854
rect 293794 329534 294414 329618
rect 293794 329298 293826 329534
rect 294062 329298 294146 329534
rect 294382 329298 294414 329534
rect 329794 329618 329826 329854
rect 330062 329618 330146 329854
rect 330382 329618 330414 329854
rect 329794 329534 330414 329618
rect 329794 329298 329826 329534
rect 330062 329298 330146 329534
rect 330382 329298 330414 329534
rect 365794 329618 365826 329854
rect 366062 329618 366146 329854
rect 366382 329618 366414 329854
rect 365794 329534 366414 329618
rect 365794 329298 365826 329534
rect 366062 329298 366146 329534
rect 366382 329298 366414 329534
rect 401794 329618 401826 329854
rect 402062 329618 402146 329854
rect 402382 329618 402414 329854
rect 401794 329534 402414 329618
rect 401794 329298 401826 329534
rect 402062 329298 402146 329534
rect 402382 329298 402414 329534
rect 570318 329618 570350 329854
rect 570586 329618 570670 329854
rect 570906 329618 570938 329854
rect 570318 329534 570938 329618
rect 570318 329298 570350 329534
rect 570586 329298 570670 329534
rect 570906 329298 570938 329534
rect -2006 293854 -1386 329298
rect 582294 298354 582914 333798
rect 13166 298118 13198 298354
rect 13434 298118 13518 298354
rect 13754 298118 13786 298354
rect 13166 298034 13786 298118
rect 13166 297798 13198 298034
rect 13434 297798 13518 298034
rect 13754 297798 13786 298034
rect 167794 298118 167826 298354
rect 168062 298118 168146 298354
rect 168382 298118 168414 298354
rect 167794 298034 168414 298118
rect 167794 297798 167826 298034
rect 168062 297798 168146 298034
rect 168382 297798 168414 298034
rect 203794 298118 203826 298354
rect 204062 298118 204146 298354
rect 204382 298118 204414 298354
rect 203794 298034 204414 298118
rect 203794 297798 203826 298034
rect 204062 297798 204146 298034
rect 204382 297798 204414 298034
rect 239794 298118 239826 298354
rect 240062 298118 240146 298354
rect 240382 298118 240414 298354
rect 239794 298034 240414 298118
rect 239794 297798 239826 298034
rect 240062 297798 240146 298034
rect 240382 297798 240414 298034
rect 275794 298118 275826 298354
rect 276062 298118 276146 298354
rect 276382 298118 276414 298354
rect 275794 298034 276414 298118
rect 275794 297798 275826 298034
rect 276062 297798 276146 298034
rect 276382 297798 276414 298034
rect 311794 298118 311826 298354
rect 312062 298118 312146 298354
rect 312382 298118 312414 298354
rect 311794 298034 312414 298118
rect 311794 297798 311826 298034
rect 312062 297798 312146 298034
rect 312382 297798 312414 298034
rect 347794 298118 347826 298354
rect 348062 298118 348146 298354
rect 348382 298118 348414 298354
rect 347794 298034 348414 298118
rect 347794 297798 347826 298034
rect 348062 297798 348146 298034
rect 348382 297798 348414 298034
rect 383794 298118 383826 298354
rect 384062 298118 384146 298354
rect 384382 298118 384414 298354
rect 383794 298034 384414 298118
rect 383794 297798 383826 298034
rect 384062 297798 384146 298034
rect 384382 297798 384414 298034
rect 419794 298118 419826 298354
rect 420062 298118 420146 298354
rect 420382 298118 420414 298354
rect 419794 298034 420414 298118
rect 419794 297798 419826 298034
rect 420062 297798 420146 298034
rect 420382 297798 420414 298034
rect 563794 298118 563826 298354
rect 564062 298118 564146 298354
rect 564382 298118 564414 298354
rect 563794 298034 564414 298118
rect 563794 297798 563826 298034
rect 564062 297798 564146 298034
rect 564382 297798 564414 298034
rect 582294 298118 582326 298354
rect 582562 298118 582646 298354
rect 582882 298118 582914 298354
rect 582294 298034 582914 298118
rect 582294 297798 582326 298034
rect 582562 297798 582646 298034
rect 582882 297798 582914 298034
rect -2006 293618 -1974 293854
rect -1738 293618 -1654 293854
rect -1418 293618 -1386 293854
rect -2006 293534 -1386 293618
rect -2006 293298 -1974 293534
rect -1738 293298 -1654 293534
rect -1418 293298 -1386 293534
rect 5794 293618 5826 293854
rect 6062 293618 6146 293854
rect 6382 293618 6414 293854
rect 5794 293534 6414 293618
rect 5794 293298 5826 293534
rect 6062 293298 6146 293534
rect 6382 293298 6414 293534
rect 185794 293618 185826 293854
rect 186062 293618 186146 293854
rect 186382 293618 186414 293854
rect 185794 293534 186414 293618
rect 185794 293298 185826 293534
rect 186062 293298 186146 293534
rect 186382 293298 186414 293534
rect 221794 293618 221826 293854
rect 222062 293618 222146 293854
rect 222382 293618 222414 293854
rect 221794 293534 222414 293618
rect 221794 293298 221826 293534
rect 222062 293298 222146 293534
rect 222382 293298 222414 293534
rect 257794 293618 257826 293854
rect 258062 293618 258146 293854
rect 258382 293618 258414 293854
rect 257794 293534 258414 293618
rect 257794 293298 257826 293534
rect 258062 293298 258146 293534
rect 258382 293298 258414 293534
rect 293794 293618 293826 293854
rect 294062 293618 294146 293854
rect 294382 293618 294414 293854
rect 293794 293534 294414 293618
rect 293794 293298 293826 293534
rect 294062 293298 294146 293534
rect 294382 293298 294414 293534
rect 329794 293618 329826 293854
rect 330062 293618 330146 293854
rect 330382 293618 330414 293854
rect 329794 293534 330414 293618
rect 329794 293298 329826 293534
rect 330062 293298 330146 293534
rect 330382 293298 330414 293534
rect 365794 293618 365826 293854
rect 366062 293618 366146 293854
rect 366382 293618 366414 293854
rect 365794 293534 366414 293618
rect 365794 293298 365826 293534
rect 366062 293298 366146 293534
rect 366382 293298 366414 293534
rect 401794 293618 401826 293854
rect 402062 293618 402146 293854
rect 402382 293618 402414 293854
rect 401794 293534 402414 293618
rect 401794 293298 401826 293534
rect 402062 293298 402146 293534
rect 402382 293298 402414 293534
rect 570318 293618 570350 293854
rect 570586 293618 570670 293854
rect 570906 293618 570938 293854
rect 570318 293534 570938 293618
rect 570318 293298 570350 293534
rect 570586 293298 570670 293534
rect 570906 293298 570938 293534
rect -2006 257854 -1386 293298
rect 582294 262354 582914 297798
rect 13166 262118 13198 262354
rect 13434 262118 13518 262354
rect 13754 262118 13786 262354
rect 13166 262034 13786 262118
rect 13166 261798 13198 262034
rect 13434 261798 13518 262034
rect 13754 261798 13786 262034
rect 167794 262118 167826 262354
rect 168062 262118 168146 262354
rect 168382 262118 168414 262354
rect 167794 262034 168414 262118
rect 167794 261798 167826 262034
rect 168062 261798 168146 262034
rect 168382 261798 168414 262034
rect 203794 262118 203826 262354
rect 204062 262118 204146 262354
rect 204382 262118 204414 262354
rect 203794 262034 204414 262118
rect 203794 261798 203826 262034
rect 204062 261798 204146 262034
rect 204382 261798 204414 262034
rect 239794 262118 239826 262354
rect 240062 262118 240146 262354
rect 240382 262118 240414 262354
rect 239794 262034 240414 262118
rect 239794 261798 239826 262034
rect 240062 261798 240146 262034
rect 240382 261798 240414 262034
rect 275794 262118 275826 262354
rect 276062 262118 276146 262354
rect 276382 262118 276414 262354
rect 275794 262034 276414 262118
rect 275794 261798 275826 262034
rect 276062 261798 276146 262034
rect 276382 261798 276414 262034
rect 311794 262118 311826 262354
rect 312062 262118 312146 262354
rect 312382 262118 312414 262354
rect 311794 262034 312414 262118
rect 311794 261798 311826 262034
rect 312062 261798 312146 262034
rect 312382 261798 312414 262034
rect 347794 262118 347826 262354
rect 348062 262118 348146 262354
rect 348382 262118 348414 262354
rect 347794 262034 348414 262118
rect 347794 261798 347826 262034
rect 348062 261798 348146 262034
rect 348382 261798 348414 262034
rect 383794 262118 383826 262354
rect 384062 262118 384146 262354
rect 384382 262118 384414 262354
rect 383794 262034 384414 262118
rect 383794 261798 383826 262034
rect 384062 261798 384146 262034
rect 384382 261798 384414 262034
rect 419794 262118 419826 262354
rect 420062 262118 420146 262354
rect 420382 262118 420414 262354
rect 419794 262034 420414 262118
rect 419794 261798 419826 262034
rect 420062 261798 420146 262034
rect 420382 261798 420414 262034
rect 563794 262118 563826 262354
rect 564062 262118 564146 262354
rect 564382 262118 564414 262354
rect 563794 262034 564414 262118
rect 563794 261798 563826 262034
rect 564062 261798 564146 262034
rect 564382 261798 564414 262034
rect 582294 262118 582326 262354
rect 582562 262118 582646 262354
rect 582882 262118 582914 262354
rect 582294 262034 582914 262118
rect 582294 261798 582326 262034
rect 582562 261798 582646 262034
rect 582882 261798 582914 262034
rect -2006 257618 -1974 257854
rect -1738 257618 -1654 257854
rect -1418 257618 -1386 257854
rect -2006 257534 -1386 257618
rect -2006 257298 -1974 257534
rect -1738 257298 -1654 257534
rect -1418 257298 -1386 257534
rect 5794 257618 5826 257854
rect 6062 257618 6146 257854
rect 6382 257618 6414 257854
rect 5794 257534 6414 257618
rect 5794 257298 5826 257534
rect 6062 257298 6146 257534
rect 6382 257298 6414 257534
rect 185794 257618 185826 257854
rect 186062 257618 186146 257854
rect 186382 257618 186414 257854
rect 185794 257534 186414 257618
rect 185794 257298 185826 257534
rect 186062 257298 186146 257534
rect 186382 257298 186414 257534
rect 221794 257618 221826 257854
rect 222062 257618 222146 257854
rect 222382 257618 222414 257854
rect 221794 257534 222414 257618
rect 221794 257298 221826 257534
rect 222062 257298 222146 257534
rect 222382 257298 222414 257534
rect 257794 257618 257826 257854
rect 258062 257618 258146 257854
rect 258382 257618 258414 257854
rect 257794 257534 258414 257618
rect 257794 257298 257826 257534
rect 258062 257298 258146 257534
rect 258382 257298 258414 257534
rect 293794 257618 293826 257854
rect 294062 257618 294146 257854
rect 294382 257618 294414 257854
rect 293794 257534 294414 257618
rect 293794 257298 293826 257534
rect 294062 257298 294146 257534
rect 294382 257298 294414 257534
rect 329794 257618 329826 257854
rect 330062 257618 330146 257854
rect 330382 257618 330414 257854
rect 329794 257534 330414 257618
rect 329794 257298 329826 257534
rect 330062 257298 330146 257534
rect 330382 257298 330414 257534
rect 365794 257618 365826 257854
rect 366062 257618 366146 257854
rect 366382 257618 366414 257854
rect 365794 257534 366414 257618
rect 365794 257298 365826 257534
rect 366062 257298 366146 257534
rect 366382 257298 366414 257534
rect 401794 257618 401826 257854
rect 402062 257618 402146 257854
rect 402382 257618 402414 257854
rect 401794 257534 402414 257618
rect 401794 257298 401826 257534
rect 402062 257298 402146 257534
rect 402382 257298 402414 257534
rect 570318 257618 570350 257854
rect 570586 257618 570670 257854
rect 570906 257618 570938 257854
rect 570318 257534 570938 257618
rect 570318 257298 570350 257534
rect 570586 257298 570670 257534
rect 570906 257298 570938 257534
rect -2006 221854 -1386 257298
rect 582294 226354 582914 261798
rect 13166 226118 13198 226354
rect 13434 226118 13518 226354
rect 13754 226118 13786 226354
rect 13166 226034 13786 226118
rect 13166 225798 13198 226034
rect 13434 225798 13518 226034
rect 13754 225798 13786 226034
rect 167794 226118 167826 226354
rect 168062 226118 168146 226354
rect 168382 226118 168414 226354
rect 167794 226034 168414 226118
rect 167794 225798 167826 226034
rect 168062 225798 168146 226034
rect 168382 225798 168414 226034
rect 203794 226118 203826 226354
rect 204062 226118 204146 226354
rect 204382 226118 204414 226354
rect 203794 226034 204414 226118
rect 203794 225798 203826 226034
rect 204062 225798 204146 226034
rect 204382 225798 204414 226034
rect 239794 226118 239826 226354
rect 240062 226118 240146 226354
rect 240382 226118 240414 226354
rect 239794 226034 240414 226118
rect 239794 225798 239826 226034
rect 240062 225798 240146 226034
rect 240382 225798 240414 226034
rect 275794 226118 275826 226354
rect 276062 226118 276146 226354
rect 276382 226118 276414 226354
rect 275794 226034 276414 226118
rect 275794 225798 275826 226034
rect 276062 225798 276146 226034
rect 276382 225798 276414 226034
rect 311794 226118 311826 226354
rect 312062 226118 312146 226354
rect 312382 226118 312414 226354
rect 311794 226034 312414 226118
rect 311794 225798 311826 226034
rect 312062 225798 312146 226034
rect 312382 225798 312414 226034
rect 347794 226118 347826 226354
rect 348062 226118 348146 226354
rect 348382 226118 348414 226354
rect 347794 226034 348414 226118
rect 347794 225798 347826 226034
rect 348062 225798 348146 226034
rect 348382 225798 348414 226034
rect 383794 226118 383826 226354
rect 384062 226118 384146 226354
rect 384382 226118 384414 226354
rect 383794 226034 384414 226118
rect 383794 225798 383826 226034
rect 384062 225798 384146 226034
rect 384382 225798 384414 226034
rect 419794 226118 419826 226354
rect 420062 226118 420146 226354
rect 420382 226118 420414 226354
rect 419794 226034 420414 226118
rect 419794 225798 419826 226034
rect 420062 225798 420146 226034
rect 420382 225798 420414 226034
rect 563794 226118 563826 226354
rect 564062 226118 564146 226354
rect 564382 226118 564414 226354
rect 563794 226034 564414 226118
rect 563794 225798 563826 226034
rect 564062 225798 564146 226034
rect 564382 225798 564414 226034
rect 582294 226118 582326 226354
rect 582562 226118 582646 226354
rect 582882 226118 582914 226354
rect 582294 226034 582914 226118
rect 582294 225798 582326 226034
rect 582562 225798 582646 226034
rect 582882 225798 582914 226034
rect -2006 221618 -1974 221854
rect -1738 221618 -1654 221854
rect -1418 221618 -1386 221854
rect -2006 221534 -1386 221618
rect -2006 221298 -1974 221534
rect -1738 221298 -1654 221534
rect -1418 221298 -1386 221534
rect 5794 221618 5826 221854
rect 6062 221618 6146 221854
rect 6382 221618 6414 221854
rect 5794 221534 6414 221618
rect 5794 221298 5826 221534
rect 6062 221298 6146 221534
rect 6382 221298 6414 221534
rect 185794 221618 185826 221854
rect 186062 221618 186146 221854
rect 186382 221618 186414 221854
rect 185794 221534 186414 221618
rect 185794 221298 185826 221534
rect 186062 221298 186146 221534
rect 186382 221298 186414 221534
rect 221794 221618 221826 221854
rect 222062 221618 222146 221854
rect 222382 221618 222414 221854
rect 221794 221534 222414 221618
rect 221794 221298 221826 221534
rect 222062 221298 222146 221534
rect 222382 221298 222414 221534
rect 257794 221618 257826 221854
rect 258062 221618 258146 221854
rect 258382 221618 258414 221854
rect 257794 221534 258414 221618
rect 257794 221298 257826 221534
rect 258062 221298 258146 221534
rect 258382 221298 258414 221534
rect 293794 221618 293826 221854
rect 294062 221618 294146 221854
rect 294382 221618 294414 221854
rect 293794 221534 294414 221618
rect 293794 221298 293826 221534
rect 294062 221298 294146 221534
rect 294382 221298 294414 221534
rect 329794 221618 329826 221854
rect 330062 221618 330146 221854
rect 330382 221618 330414 221854
rect 329794 221534 330414 221618
rect 329794 221298 329826 221534
rect 330062 221298 330146 221534
rect 330382 221298 330414 221534
rect 365794 221618 365826 221854
rect 366062 221618 366146 221854
rect 366382 221618 366414 221854
rect 365794 221534 366414 221618
rect 365794 221298 365826 221534
rect 366062 221298 366146 221534
rect 366382 221298 366414 221534
rect 401794 221618 401826 221854
rect 402062 221618 402146 221854
rect 402382 221618 402414 221854
rect 401794 221534 402414 221618
rect 401794 221298 401826 221534
rect 402062 221298 402146 221534
rect 402382 221298 402414 221534
rect 570318 221618 570350 221854
rect 570586 221618 570670 221854
rect 570906 221618 570938 221854
rect 570318 221534 570938 221618
rect 570318 221298 570350 221534
rect 570586 221298 570670 221534
rect 570906 221298 570938 221534
rect -2006 185854 -1386 221298
rect 582294 190354 582914 225798
rect 13166 190118 13198 190354
rect 13434 190118 13518 190354
rect 13754 190118 13786 190354
rect 13166 190034 13786 190118
rect 13166 189798 13198 190034
rect 13434 189798 13518 190034
rect 13754 189798 13786 190034
rect 167794 190118 167826 190354
rect 168062 190118 168146 190354
rect 168382 190118 168414 190354
rect 167794 190034 168414 190118
rect 167794 189798 167826 190034
rect 168062 189798 168146 190034
rect 168382 189798 168414 190034
rect 203794 190118 203826 190354
rect 204062 190118 204146 190354
rect 204382 190118 204414 190354
rect 203794 190034 204414 190118
rect 203794 189798 203826 190034
rect 204062 189798 204146 190034
rect 204382 189798 204414 190034
rect 239794 190118 239826 190354
rect 240062 190118 240146 190354
rect 240382 190118 240414 190354
rect 239794 190034 240414 190118
rect 239794 189798 239826 190034
rect 240062 189798 240146 190034
rect 240382 189798 240414 190034
rect 275794 190118 275826 190354
rect 276062 190118 276146 190354
rect 276382 190118 276414 190354
rect 275794 190034 276414 190118
rect 275794 189798 275826 190034
rect 276062 189798 276146 190034
rect 276382 189798 276414 190034
rect 311794 190118 311826 190354
rect 312062 190118 312146 190354
rect 312382 190118 312414 190354
rect 311794 190034 312414 190118
rect 311794 189798 311826 190034
rect 312062 189798 312146 190034
rect 312382 189798 312414 190034
rect 347794 190118 347826 190354
rect 348062 190118 348146 190354
rect 348382 190118 348414 190354
rect 347794 190034 348414 190118
rect 347794 189798 347826 190034
rect 348062 189798 348146 190034
rect 348382 189798 348414 190034
rect 383794 190118 383826 190354
rect 384062 190118 384146 190354
rect 384382 190118 384414 190354
rect 383794 190034 384414 190118
rect 383794 189798 383826 190034
rect 384062 189798 384146 190034
rect 384382 189798 384414 190034
rect 419794 190118 419826 190354
rect 420062 190118 420146 190354
rect 420382 190118 420414 190354
rect 419794 190034 420414 190118
rect 419794 189798 419826 190034
rect 420062 189798 420146 190034
rect 420382 189798 420414 190034
rect 563794 190118 563826 190354
rect 564062 190118 564146 190354
rect 564382 190118 564414 190354
rect 563794 190034 564414 190118
rect 563794 189798 563826 190034
rect 564062 189798 564146 190034
rect 564382 189798 564414 190034
rect 582294 190118 582326 190354
rect 582562 190118 582646 190354
rect 582882 190118 582914 190354
rect 582294 190034 582914 190118
rect 582294 189798 582326 190034
rect 582562 189798 582646 190034
rect 582882 189798 582914 190034
rect -2006 185618 -1974 185854
rect -1738 185618 -1654 185854
rect -1418 185618 -1386 185854
rect -2006 185534 -1386 185618
rect -2006 185298 -1974 185534
rect -1738 185298 -1654 185534
rect -1418 185298 -1386 185534
rect 5794 185618 5826 185854
rect 6062 185618 6146 185854
rect 6382 185618 6414 185854
rect 5794 185534 6414 185618
rect 5794 185298 5826 185534
rect 6062 185298 6146 185534
rect 6382 185298 6414 185534
rect 185794 185618 185826 185854
rect 186062 185618 186146 185854
rect 186382 185618 186414 185854
rect 185794 185534 186414 185618
rect 185794 185298 185826 185534
rect 186062 185298 186146 185534
rect 186382 185298 186414 185534
rect 221794 185618 221826 185854
rect 222062 185618 222146 185854
rect 222382 185618 222414 185854
rect 221794 185534 222414 185618
rect 221794 185298 221826 185534
rect 222062 185298 222146 185534
rect 222382 185298 222414 185534
rect 257794 185618 257826 185854
rect 258062 185618 258146 185854
rect 258382 185618 258414 185854
rect 257794 185534 258414 185618
rect 257794 185298 257826 185534
rect 258062 185298 258146 185534
rect 258382 185298 258414 185534
rect 293794 185618 293826 185854
rect 294062 185618 294146 185854
rect 294382 185618 294414 185854
rect 293794 185534 294414 185618
rect 293794 185298 293826 185534
rect 294062 185298 294146 185534
rect 294382 185298 294414 185534
rect 329794 185618 329826 185854
rect 330062 185618 330146 185854
rect 330382 185618 330414 185854
rect 329794 185534 330414 185618
rect 329794 185298 329826 185534
rect 330062 185298 330146 185534
rect 330382 185298 330414 185534
rect 365794 185618 365826 185854
rect 366062 185618 366146 185854
rect 366382 185618 366414 185854
rect 365794 185534 366414 185618
rect 365794 185298 365826 185534
rect 366062 185298 366146 185534
rect 366382 185298 366414 185534
rect 401794 185618 401826 185854
rect 402062 185618 402146 185854
rect 402382 185618 402414 185854
rect 401794 185534 402414 185618
rect 401794 185298 401826 185534
rect 402062 185298 402146 185534
rect 402382 185298 402414 185534
rect 570318 185618 570350 185854
rect 570586 185618 570670 185854
rect 570906 185618 570938 185854
rect 570318 185534 570938 185618
rect 570318 185298 570350 185534
rect 570586 185298 570670 185534
rect 570906 185298 570938 185534
rect -2006 149854 -1386 185298
rect 582294 154354 582914 189798
rect 13166 154118 13198 154354
rect 13434 154118 13518 154354
rect 13754 154118 13786 154354
rect 13166 154034 13786 154118
rect 13166 153798 13198 154034
rect 13434 153798 13518 154034
rect 13754 153798 13786 154034
rect 167794 154118 167826 154354
rect 168062 154118 168146 154354
rect 168382 154118 168414 154354
rect 167794 154034 168414 154118
rect 167794 153798 167826 154034
rect 168062 153798 168146 154034
rect 168382 153798 168414 154034
rect 203794 154118 203826 154354
rect 204062 154118 204146 154354
rect 204382 154118 204414 154354
rect 203794 154034 204414 154118
rect 203794 153798 203826 154034
rect 204062 153798 204146 154034
rect 204382 153798 204414 154034
rect 239794 154118 239826 154354
rect 240062 154118 240146 154354
rect 240382 154118 240414 154354
rect 239794 154034 240414 154118
rect 239794 153798 239826 154034
rect 240062 153798 240146 154034
rect 240382 153798 240414 154034
rect 275794 154118 275826 154354
rect 276062 154118 276146 154354
rect 276382 154118 276414 154354
rect 275794 154034 276414 154118
rect 275794 153798 275826 154034
rect 276062 153798 276146 154034
rect 276382 153798 276414 154034
rect 311794 154118 311826 154354
rect 312062 154118 312146 154354
rect 312382 154118 312414 154354
rect 311794 154034 312414 154118
rect 311794 153798 311826 154034
rect 312062 153798 312146 154034
rect 312382 153798 312414 154034
rect 347794 154118 347826 154354
rect 348062 154118 348146 154354
rect 348382 154118 348414 154354
rect 347794 154034 348414 154118
rect 347794 153798 347826 154034
rect 348062 153798 348146 154034
rect 348382 153798 348414 154034
rect 383794 154118 383826 154354
rect 384062 154118 384146 154354
rect 384382 154118 384414 154354
rect 383794 154034 384414 154118
rect 383794 153798 383826 154034
rect 384062 153798 384146 154034
rect 384382 153798 384414 154034
rect 419794 154118 419826 154354
rect 420062 154118 420146 154354
rect 420382 154118 420414 154354
rect 419794 154034 420414 154118
rect 419794 153798 419826 154034
rect 420062 153798 420146 154034
rect 420382 153798 420414 154034
rect 563794 154118 563826 154354
rect 564062 154118 564146 154354
rect 564382 154118 564414 154354
rect 563794 154034 564414 154118
rect 563794 153798 563826 154034
rect 564062 153798 564146 154034
rect 564382 153798 564414 154034
rect 582294 154118 582326 154354
rect 582562 154118 582646 154354
rect 582882 154118 582914 154354
rect 582294 154034 582914 154118
rect 582294 153798 582326 154034
rect 582562 153798 582646 154034
rect 582882 153798 582914 154034
rect -2006 149618 -1974 149854
rect -1738 149618 -1654 149854
rect -1418 149618 -1386 149854
rect -2006 149534 -1386 149618
rect -2006 149298 -1974 149534
rect -1738 149298 -1654 149534
rect -1418 149298 -1386 149534
rect 5794 149618 5826 149854
rect 6062 149618 6146 149854
rect 6382 149618 6414 149854
rect 5794 149534 6414 149618
rect 5794 149298 5826 149534
rect 6062 149298 6146 149534
rect 6382 149298 6414 149534
rect 185794 149618 185826 149854
rect 186062 149618 186146 149854
rect 186382 149618 186414 149854
rect 185794 149534 186414 149618
rect 185794 149298 185826 149534
rect 186062 149298 186146 149534
rect 186382 149298 186414 149534
rect 221794 149618 221826 149854
rect 222062 149618 222146 149854
rect 222382 149618 222414 149854
rect 221794 149534 222414 149618
rect 221794 149298 221826 149534
rect 222062 149298 222146 149534
rect 222382 149298 222414 149534
rect 257794 149618 257826 149854
rect 258062 149618 258146 149854
rect 258382 149618 258414 149854
rect 257794 149534 258414 149618
rect 257794 149298 257826 149534
rect 258062 149298 258146 149534
rect 258382 149298 258414 149534
rect 293794 149618 293826 149854
rect 294062 149618 294146 149854
rect 294382 149618 294414 149854
rect 293794 149534 294414 149618
rect 293794 149298 293826 149534
rect 294062 149298 294146 149534
rect 294382 149298 294414 149534
rect 329794 149618 329826 149854
rect 330062 149618 330146 149854
rect 330382 149618 330414 149854
rect 329794 149534 330414 149618
rect 329794 149298 329826 149534
rect 330062 149298 330146 149534
rect 330382 149298 330414 149534
rect 365794 149618 365826 149854
rect 366062 149618 366146 149854
rect 366382 149618 366414 149854
rect 365794 149534 366414 149618
rect 365794 149298 365826 149534
rect 366062 149298 366146 149534
rect 366382 149298 366414 149534
rect 401794 149618 401826 149854
rect 402062 149618 402146 149854
rect 402382 149618 402414 149854
rect 401794 149534 402414 149618
rect 401794 149298 401826 149534
rect 402062 149298 402146 149534
rect 402382 149298 402414 149534
rect 570318 149618 570350 149854
rect 570586 149618 570670 149854
rect 570906 149618 570938 149854
rect 570318 149534 570938 149618
rect 570318 149298 570350 149534
rect 570586 149298 570670 149534
rect 570906 149298 570938 149534
rect -2006 113854 -1386 149298
rect 582294 118354 582914 153798
rect 13166 118118 13198 118354
rect 13434 118118 13518 118354
rect 13754 118118 13786 118354
rect 13166 118034 13786 118118
rect 13166 117798 13198 118034
rect 13434 117798 13518 118034
rect 13754 117798 13786 118034
rect 167794 118118 167826 118354
rect 168062 118118 168146 118354
rect 168382 118118 168414 118354
rect 167794 118034 168414 118118
rect 167794 117798 167826 118034
rect 168062 117798 168146 118034
rect 168382 117798 168414 118034
rect 203794 118118 203826 118354
rect 204062 118118 204146 118354
rect 204382 118118 204414 118354
rect 203794 118034 204414 118118
rect 203794 117798 203826 118034
rect 204062 117798 204146 118034
rect 204382 117798 204414 118034
rect 239794 118118 239826 118354
rect 240062 118118 240146 118354
rect 240382 118118 240414 118354
rect 239794 118034 240414 118118
rect 239794 117798 239826 118034
rect 240062 117798 240146 118034
rect 240382 117798 240414 118034
rect 275794 118118 275826 118354
rect 276062 118118 276146 118354
rect 276382 118118 276414 118354
rect 275794 118034 276414 118118
rect 275794 117798 275826 118034
rect 276062 117798 276146 118034
rect 276382 117798 276414 118034
rect 311794 118118 311826 118354
rect 312062 118118 312146 118354
rect 312382 118118 312414 118354
rect 311794 118034 312414 118118
rect 311794 117798 311826 118034
rect 312062 117798 312146 118034
rect 312382 117798 312414 118034
rect 347794 118118 347826 118354
rect 348062 118118 348146 118354
rect 348382 118118 348414 118354
rect 347794 118034 348414 118118
rect 347794 117798 347826 118034
rect 348062 117798 348146 118034
rect 348382 117798 348414 118034
rect 383794 118118 383826 118354
rect 384062 118118 384146 118354
rect 384382 118118 384414 118354
rect 383794 118034 384414 118118
rect 383794 117798 383826 118034
rect 384062 117798 384146 118034
rect 384382 117798 384414 118034
rect 419794 118118 419826 118354
rect 420062 118118 420146 118354
rect 420382 118118 420414 118354
rect 419794 118034 420414 118118
rect 419794 117798 419826 118034
rect 420062 117798 420146 118034
rect 420382 117798 420414 118034
rect 563794 118118 563826 118354
rect 564062 118118 564146 118354
rect 564382 118118 564414 118354
rect 563794 118034 564414 118118
rect 563794 117798 563826 118034
rect 564062 117798 564146 118034
rect 564382 117798 564414 118034
rect 582294 118118 582326 118354
rect 582562 118118 582646 118354
rect 582882 118118 582914 118354
rect 582294 118034 582914 118118
rect 582294 117798 582326 118034
rect 582562 117798 582646 118034
rect 582882 117798 582914 118034
rect -2006 113618 -1974 113854
rect -1738 113618 -1654 113854
rect -1418 113618 -1386 113854
rect -2006 113534 -1386 113618
rect -2006 113298 -1974 113534
rect -1738 113298 -1654 113534
rect -1418 113298 -1386 113534
rect 5794 113618 5826 113854
rect 6062 113618 6146 113854
rect 6382 113618 6414 113854
rect 5794 113534 6414 113618
rect 5794 113298 5826 113534
rect 6062 113298 6146 113534
rect 6382 113298 6414 113534
rect 173062 113618 173094 113854
rect 173330 113618 173414 113854
rect 173650 113618 173682 113854
rect 173062 113534 173682 113618
rect 173062 113298 173094 113534
rect 173330 113298 173414 113534
rect 173650 113298 173682 113534
rect 293794 113618 293826 113854
rect 294062 113618 294146 113854
rect 294382 113618 294414 113854
rect 293794 113534 294414 113618
rect 293794 113298 293826 113534
rect 294062 113298 294146 113534
rect 294382 113298 294414 113534
rect 401794 113618 401826 113854
rect 402062 113618 402146 113854
rect 402382 113618 402414 113854
rect 401794 113534 402414 113618
rect 401794 113298 401826 113534
rect 402062 113298 402146 113534
rect 402382 113298 402414 113534
rect 570318 113618 570350 113854
rect 570586 113618 570670 113854
rect 570906 113618 570938 113854
rect 570318 113534 570938 113618
rect 570318 113298 570350 113534
rect 570586 113298 570670 113534
rect 570906 113298 570938 113534
rect -2006 77854 -1386 113298
rect 582294 82354 582914 117798
rect 13166 82118 13198 82354
rect 13434 82118 13518 82354
rect 13754 82118 13786 82354
rect 13166 82034 13786 82118
rect 13166 81798 13198 82034
rect 13434 81798 13518 82034
rect 13754 81798 13786 82034
rect 167794 82118 167826 82354
rect 168062 82118 168146 82354
rect 168382 82118 168414 82354
rect 167794 82034 168414 82118
rect 167794 81798 167826 82034
rect 168062 81798 168146 82034
rect 168382 81798 168414 82034
rect 291558 82118 291590 82354
rect 291826 82118 291910 82354
rect 292146 82118 292178 82354
rect 291558 82034 292178 82118
rect 291558 81798 291590 82034
rect 291826 81798 291910 82034
rect 292146 81798 292178 82034
rect 419794 82118 419826 82354
rect 420062 82118 420146 82354
rect 420382 82118 420414 82354
rect 419794 82034 420414 82118
rect 419794 81798 419826 82034
rect 420062 81798 420146 82034
rect 420382 81798 420414 82034
rect 563794 82118 563826 82354
rect 564062 82118 564146 82354
rect 564382 82118 564414 82354
rect 563794 82034 564414 82118
rect 563794 81798 563826 82034
rect 564062 81798 564146 82034
rect 564382 81798 564414 82034
rect 582294 82118 582326 82354
rect 582562 82118 582646 82354
rect 582882 82118 582914 82354
rect 582294 82034 582914 82118
rect 582294 81798 582326 82034
rect 582562 81798 582646 82034
rect 582882 81798 582914 82034
rect -2006 77618 -1974 77854
rect -1738 77618 -1654 77854
rect -1418 77618 -1386 77854
rect -2006 77534 -1386 77618
rect -2006 77298 -1974 77534
rect -1738 77298 -1654 77534
rect -1418 77298 -1386 77534
rect 5794 77618 5826 77854
rect 6062 77618 6146 77854
rect 6382 77618 6414 77854
rect 5794 77534 6414 77618
rect 5794 77298 5826 77534
rect 6062 77298 6146 77534
rect 6382 77298 6414 77534
rect 173062 77618 173094 77854
rect 173330 77618 173414 77854
rect 173650 77618 173682 77854
rect 173062 77534 173682 77618
rect 173062 77298 173094 77534
rect 173330 77298 173414 77534
rect 173650 77298 173682 77534
rect 293794 77618 293826 77854
rect 294062 77618 294146 77854
rect 294382 77618 294414 77854
rect 293794 77534 294414 77618
rect 293794 77298 293826 77534
rect 294062 77298 294146 77534
rect 294382 77298 294414 77534
rect 401794 77618 401826 77854
rect 402062 77618 402146 77854
rect 402382 77618 402414 77854
rect 401794 77534 402414 77618
rect 401794 77298 401826 77534
rect 402062 77298 402146 77534
rect 402382 77298 402414 77534
rect 570318 77618 570350 77854
rect 570586 77618 570670 77854
rect 570906 77618 570938 77854
rect 570318 77534 570938 77618
rect 570318 77298 570350 77534
rect 570586 77298 570670 77534
rect 570906 77298 570938 77534
rect -2006 41854 -1386 77298
rect 582294 46354 582914 81798
rect 13166 46118 13198 46354
rect 13434 46118 13518 46354
rect 13754 46118 13786 46354
rect 13166 46034 13786 46118
rect 13166 45798 13198 46034
rect 13434 45798 13518 46034
rect 13754 45798 13786 46034
rect 167794 46118 167826 46354
rect 168062 46118 168146 46354
rect 168382 46118 168414 46354
rect 167794 46034 168414 46118
rect 167794 45798 167826 46034
rect 168062 45798 168146 46034
rect 168382 45798 168414 46034
rect 291558 46118 291590 46354
rect 291826 46118 291910 46354
rect 292146 46118 292178 46354
rect 291558 46034 292178 46118
rect 291558 45798 291590 46034
rect 291826 45798 291910 46034
rect 292146 45798 292178 46034
rect 419794 46118 419826 46354
rect 420062 46118 420146 46354
rect 420382 46118 420414 46354
rect 419794 46034 420414 46118
rect 419794 45798 419826 46034
rect 420062 45798 420146 46034
rect 420382 45798 420414 46034
rect 563794 46118 563826 46354
rect 564062 46118 564146 46354
rect 564382 46118 564414 46354
rect 563794 46034 564414 46118
rect 563794 45798 563826 46034
rect 564062 45798 564146 46034
rect 564382 45798 564414 46034
rect 582294 46118 582326 46354
rect 582562 46118 582646 46354
rect 582882 46118 582914 46354
rect 582294 46034 582914 46118
rect 582294 45798 582326 46034
rect 582562 45798 582646 46034
rect 582882 45798 582914 46034
rect -2006 41618 -1974 41854
rect -1738 41618 -1654 41854
rect -1418 41618 -1386 41854
rect -2006 41534 -1386 41618
rect -2006 41298 -1974 41534
rect -1738 41298 -1654 41534
rect -1418 41298 -1386 41534
rect 5794 41618 5826 41854
rect 6062 41618 6146 41854
rect 6382 41618 6414 41854
rect 5794 41534 6414 41618
rect 5794 41298 5826 41534
rect 6062 41298 6146 41534
rect 6382 41298 6414 41534
rect 173062 41618 173094 41854
rect 173330 41618 173414 41854
rect 173650 41618 173682 41854
rect 173062 41534 173682 41618
rect 173062 41298 173094 41534
rect 173330 41298 173414 41534
rect 173650 41298 173682 41534
rect 293794 41618 293826 41854
rect 294062 41618 294146 41854
rect 294382 41618 294414 41854
rect 293794 41534 294414 41618
rect 293794 41298 293826 41534
rect 294062 41298 294146 41534
rect 294382 41298 294414 41534
rect 401794 41618 401826 41854
rect 402062 41618 402146 41854
rect 402382 41618 402414 41854
rect 401794 41534 402414 41618
rect 401794 41298 401826 41534
rect 402062 41298 402146 41534
rect 402382 41298 402414 41534
rect 570318 41618 570350 41854
rect 570586 41618 570670 41854
rect 570906 41618 570938 41854
rect 570318 41534 570938 41618
rect 570318 41298 570350 41534
rect 570586 41298 570670 41534
rect 570906 41298 570938 41534
rect -2006 5854 -1386 41298
rect 582294 10354 582914 45798
rect 23794 10118 23826 10354
rect 24062 10118 24146 10354
rect 24382 10118 24414 10354
rect 23794 10034 24414 10118
rect 23794 9798 23826 10034
rect 24062 9798 24146 10034
rect 24382 9798 24414 10034
rect 59794 10118 59826 10354
rect 60062 10118 60146 10354
rect 60382 10118 60414 10354
rect 59794 10034 60414 10118
rect 59794 9798 59826 10034
rect 60062 9798 60146 10034
rect 60382 9798 60414 10034
rect 95794 10118 95826 10354
rect 96062 10118 96146 10354
rect 96382 10118 96414 10354
rect 95794 10034 96414 10118
rect 95794 9798 95826 10034
rect 96062 9798 96146 10034
rect 96382 9798 96414 10034
rect 131794 10118 131826 10354
rect 132062 10118 132146 10354
rect 132382 10118 132414 10354
rect 131794 10034 132414 10118
rect 131794 9798 131826 10034
rect 132062 9798 132146 10034
rect 132382 9798 132414 10034
rect 167794 10118 167826 10354
rect 168062 10118 168146 10354
rect 168382 10118 168414 10354
rect 167794 10034 168414 10118
rect 167794 9798 167826 10034
rect 168062 9798 168146 10034
rect 168382 9798 168414 10034
rect 203794 10118 203826 10354
rect 204062 10118 204146 10354
rect 204382 10118 204414 10354
rect 203794 10034 204414 10118
rect 203794 9798 203826 10034
rect 204062 9798 204146 10034
rect 204382 9798 204414 10034
rect 239794 10118 239826 10354
rect 240062 10118 240146 10354
rect 240382 10118 240414 10354
rect 239794 10034 240414 10118
rect 239794 9798 239826 10034
rect 240062 9798 240146 10034
rect 240382 9798 240414 10034
rect 275794 10118 275826 10354
rect 276062 10118 276146 10354
rect 276382 10118 276414 10354
rect 275794 10034 276414 10118
rect 275794 9798 275826 10034
rect 276062 9798 276146 10034
rect 276382 9798 276414 10034
rect 311794 10118 311826 10354
rect 312062 10118 312146 10354
rect 312382 10118 312414 10354
rect 311794 10034 312414 10118
rect 311794 9798 311826 10034
rect 312062 9798 312146 10034
rect 312382 9798 312414 10034
rect 347794 10118 347826 10354
rect 348062 10118 348146 10354
rect 348382 10118 348414 10354
rect 347794 10034 348414 10118
rect 347794 9798 347826 10034
rect 348062 9798 348146 10034
rect 348382 9798 348414 10034
rect 383794 10118 383826 10354
rect 384062 10118 384146 10354
rect 384382 10118 384414 10354
rect 383794 10034 384414 10118
rect 383794 9798 383826 10034
rect 384062 9798 384146 10034
rect 384382 9798 384414 10034
rect 419794 10118 419826 10354
rect 420062 10118 420146 10354
rect 420382 10118 420414 10354
rect 419794 10034 420414 10118
rect 419794 9798 419826 10034
rect 420062 9798 420146 10034
rect 420382 9798 420414 10034
rect 455794 10118 455826 10354
rect 456062 10118 456146 10354
rect 456382 10118 456414 10354
rect 455794 10034 456414 10118
rect 455794 9798 455826 10034
rect 456062 9798 456146 10034
rect 456382 9798 456414 10034
rect 491794 10118 491826 10354
rect 492062 10118 492146 10354
rect 492382 10118 492414 10354
rect 491794 10034 492414 10118
rect 491794 9798 491826 10034
rect 492062 9798 492146 10034
rect 492382 9798 492414 10034
rect 527794 10118 527826 10354
rect 528062 10118 528146 10354
rect 528382 10118 528414 10354
rect 527794 10034 528414 10118
rect 527794 9798 527826 10034
rect 528062 9798 528146 10034
rect 528382 9798 528414 10034
rect 563794 10118 563826 10354
rect 564062 10118 564146 10354
rect 564382 10118 564414 10354
rect 563794 10034 564414 10118
rect 563794 9798 563826 10034
rect 564062 9798 564146 10034
rect 564382 9798 564414 10034
rect 582294 10118 582326 10354
rect 582562 10118 582646 10354
rect 582882 10118 582914 10354
rect 582294 10034 582914 10118
rect 582294 9798 582326 10034
rect 582562 9798 582646 10034
rect 582882 9798 582914 10034
rect -2006 5618 -1974 5854
rect -1738 5618 -1654 5854
rect -1418 5618 -1386 5854
rect -2006 5534 -1386 5618
rect -2006 5298 -1974 5534
rect -1738 5298 -1654 5534
rect -1418 5298 -1386 5534
rect -2006 -346 -1386 5298
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect 582294 -1306 582914 9798
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 689854 585930 704282
rect 585310 689618 585342 689854
rect 585578 689618 585662 689854
rect 585898 689618 585930 689854
rect 585310 689534 585930 689618
rect 585310 689298 585342 689534
rect 585578 689298 585662 689534
rect 585898 689298 585930 689534
rect 585310 653854 585930 689298
rect 585310 653618 585342 653854
rect 585578 653618 585662 653854
rect 585898 653618 585930 653854
rect 585310 653534 585930 653618
rect 585310 653298 585342 653534
rect 585578 653298 585662 653534
rect 585898 653298 585930 653534
rect 585310 617854 585930 653298
rect 585310 617618 585342 617854
rect 585578 617618 585662 617854
rect 585898 617618 585930 617854
rect 585310 617534 585930 617618
rect 585310 617298 585342 617534
rect 585578 617298 585662 617534
rect 585898 617298 585930 617534
rect 585310 581854 585930 617298
rect 585310 581618 585342 581854
rect 585578 581618 585662 581854
rect 585898 581618 585930 581854
rect 585310 581534 585930 581618
rect 585310 581298 585342 581534
rect 585578 581298 585662 581534
rect 585898 581298 585930 581534
rect 585310 545854 585930 581298
rect 585310 545618 585342 545854
rect 585578 545618 585662 545854
rect 585898 545618 585930 545854
rect 585310 545534 585930 545618
rect 585310 545298 585342 545534
rect 585578 545298 585662 545534
rect 585898 545298 585930 545534
rect 585310 509854 585930 545298
rect 585310 509618 585342 509854
rect 585578 509618 585662 509854
rect 585898 509618 585930 509854
rect 585310 509534 585930 509618
rect 585310 509298 585342 509534
rect 585578 509298 585662 509534
rect 585898 509298 585930 509534
rect 585310 473854 585930 509298
rect 585310 473618 585342 473854
rect 585578 473618 585662 473854
rect 585898 473618 585930 473854
rect 585310 473534 585930 473618
rect 585310 473298 585342 473534
rect 585578 473298 585662 473534
rect 585898 473298 585930 473534
rect 585310 437854 585930 473298
rect 585310 437618 585342 437854
rect 585578 437618 585662 437854
rect 585898 437618 585930 437854
rect 585310 437534 585930 437618
rect 585310 437298 585342 437534
rect 585578 437298 585662 437534
rect 585898 437298 585930 437534
rect 585310 401854 585930 437298
rect 585310 401618 585342 401854
rect 585578 401618 585662 401854
rect 585898 401618 585930 401854
rect 585310 401534 585930 401618
rect 585310 401298 585342 401534
rect 585578 401298 585662 401534
rect 585898 401298 585930 401534
rect 585310 365854 585930 401298
rect 585310 365618 585342 365854
rect 585578 365618 585662 365854
rect 585898 365618 585930 365854
rect 585310 365534 585930 365618
rect 585310 365298 585342 365534
rect 585578 365298 585662 365534
rect 585898 365298 585930 365534
rect 585310 329854 585930 365298
rect 585310 329618 585342 329854
rect 585578 329618 585662 329854
rect 585898 329618 585930 329854
rect 585310 329534 585930 329618
rect 585310 329298 585342 329534
rect 585578 329298 585662 329534
rect 585898 329298 585930 329534
rect 585310 293854 585930 329298
rect 585310 293618 585342 293854
rect 585578 293618 585662 293854
rect 585898 293618 585930 293854
rect 585310 293534 585930 293618
rect 585310 293298 585342 293534
rect 585578 293298 585662 293534
rect 585898 293298 585930 293534
rect 585310 257854 585930 293298
rect 585310 257618 585342 257854
rect 585578 257618 585662 257854
rect 585898 257618 585930 257854
rect 585310 257534 585930 257618
rect 585310 257298 585342 257534
rect 585578 257298 585662 257534
rect 585898 257298 585930 257534
rect 585310 221854 585930 257298
rect 585310 221618 585342 221854
rect 585578 221618 585662 221854
rect 585898 221618 585930 221854
rect 585310 221534 585930 221618
rect 585310 221298 585342 221534
rect 585578 221298 585662 221534
rect 585898 221298 585930 221534
rect 585310 185854 585930 221298
rect 585310 185618 585342 185854
rect 585578 185618 585662 185854
rect 585898 185618 585930 185854
rect 585310 185534 585930 185618
rect 585310 185298 585342 185534
rect 585578 185298 585662 185534
rect 585898 185298 585930 185534
rect 585310 149854 585930 185298
rect 585310 149618 585342 149854
rect 585578 149618 585662 149854
rect 585898 149618 585930 149854
rect 585310 149534 585930 149618
rect 585310 149298 585342 149534
rect 585578 149298 585662 149534
rect 585898 149298 585930 149534
rect 585310 113854 585930 149298
rect 585310 113618 585342 113854
rect 585578 113618 585662 113854
rect 585898 113618 585930 113854
rect 585310 113534 585930 113618
rect 585310 113298 585342 113534
rect 585578 113298 585662 113534
rect 585898 113298 585930 113534
rect 585310 77854 585930 113298
rect 585310 77618 585342 77854
rect 585578 77618 585662 77854
rect 585898 77618 585930 77854
rect 585310 77534 585930 77618
rect 585310 77298 585342 77534
rect 585578 77298 585662 77534
rect 585898 77298 585930 77534
rect 585310 41854 585930 77298
rect 585310 41618 585342 41854
rect 585578 41618 585662 41854
rect 585898 41618 585930 41854
rect 585310 41534 585930 41618
rect 585310 41298 585342 41534
rect 585578 41298 585662 41534
rect 585898 41298 585930 41534
rect 585310 5854 585930 41298
rect 585310 5618 585342 5854
rect 585578 5618 585662 5854
rect 585898 5618 585930 5854
rect 585310 5534 585930 5618
rect 585310 5298 585342 5534
rect 585578 5298 585662 5534
rect 585898 5298 585930 5534
rect 585310 -346 585930 5298
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 694354 586890 705242
rect 586270 694118 586302 694354
rect 586538 694118 586622 694354
rect 586858 694118 586890 694354
rect 586270 694034 586890 694118
rect 586270 693798 586302 694034
rect 586538 693798 586622 694034
rect 586858 693798 586890 694034
rect 586270 658354 586890 693798
rect 586270 658118 586302 658354
rect 586538 658118 586622 658354
rect 586858 658118 586890 658354
rect 586270 658034 586890 658118
rect 586270 657798 586302 658034
rect 586538 657798 586622 658034
rect 586858 657798 586890 658034
rect 586270 622354 586890 657798
rect 586270 622118 586302 622354
rect 586538 622118 586622 622354
rect 586858 622118 586890 622354
rect 586270 622034 586890 622118
rect 586270 621798 586302 622034
rect 586538 621798 586622 622034
rect 586858 621798 586890 622034
rect 586270 586354 586890 621798
rect 586270 586118 586302 586354
rect 586538 586118 586622 586354
rect 586858 586118 586890 586354
rect 586270 586034 586890 586118
rect 586270 585798 586302 586034
rect 586538 585798 586622 586034
rect 586858 585798 586890 586034
rect 586270 550354 586890 585798
rect 586270 550118 586302 550354
rect 586538 550118 586622 550354
rect 586858 550118 586890 550354
rect 586270 550034 586890 550118
rect 586270 549798 586302 550034
rect 586538 549798 586622 550034
rect 586858 549798 586890 550034
rect 586270 514354 586890 549798
rect 586270 514118 586302 514354
rect 586538 514118 586622 514354
rect 586858 514118 586890 514354
rect 586270 514034 586890 514118
rect 586270 513798 586302 514034
rect 586538 513798 586622 514034
rect 586858 513798 586890 514034
rect 586270 478354 586890 513798
rect 586270 478118 586302 478354
rect 586538 478118 586622 478354
rect 586858 478118 586890 478354
rect 586270 478034 586890 478118
rect 586270 477798 586302 478034
rect 586538 477798 586622 478034
rect 586858 477798 586890 478034
rect 586270 442354 586890 477798
rect 586270 442118 586302 442354
rect 586538 442118 586622 442354
rect 586858 442118 586890 442354
rect 586270 442034 586890 442118
rect 586270 441798 586302 442034
rect 586538 441798 586622 442034
rect 586858 441798 586890 442034
rect 586270 406354 586890 441798
rect 586270 406118 586302 406354
rect 586538 406118 586622 406354
rect 586858 406118 586890 406354
rect 586270 406034 586890 406118
rect 586270 405798 586302 406034
rect 586538 405798 586622 406034
rect 586858 405798 586890 406034
rect 586270 370354 586890 405798
rect 586270 370118 586302 370354
rect 586538 370118 586622 370354
rect 586858 370118 586890 370354
rect 586270 370034 586890 370118
rect 586270 369798 586302 370034
rect 586538 369798 586622 370034
rect 586858 369798 586890 370034
rect 586270 334354 586890 369798
rect 586270 334118 586302 334354
rect 586538 334118 586622 334354
rect 586858 334118 586890 334354
rect 586270 334034 586890 334118
rect 586270 333798 586302 334034
rect 586538 333798 586622 334034
rect 586858 333798 586890 334034
rect 586270 298354 586890 333798
rect 586270 298118 586302 298354
rect 586538 298118 586622 298354
rect 586858 298118 586890 298354
rect 586270 298034 586890 298118
rect 586270 297798 586302 298034
rect 586538 297798 586622 298034
rect 586858 297798 586890 298034
rect 586270 262354 586890 297798
rect 586270 262118 586302 262354
rect 586538 262118 586622 262354
rect 586858 262118 586890 262354
rect 586270 262034 586890 262118
rect 586270 261798 586302 262034
rect 586538 261798 586622 262034
rect 586858 261798 586890 262034
rect 586270 226354 586890 261798
rect 586270 226118 586302 226354
rect 586538 226118 586622 226354
rect 586858 226118 586890 226354
rect 586270 226034 586890 226118
rect 586270 225798 586302 226034
rect 586538 225798 586622 226034
rect 586858 225798 586890 226034
rect 586270 190354 586890 225798
rect 586270 190118 586302 190354
rect 586538 190118 586622 190354
rect 586858 190118 586890 190354
rect 586270 190034 586890 190118
rect 586270 189798 586302 190034
rect 586538 189798 586622 190034
rect 586858 189798 586890 190034
rect 586270 154354 586890 189798
rect 586270 154118 586302 154354
rect 586538 154118 586622 154354
rect 586858 154118 586890 154354
rect 586270 154034 586890 154118
rect 586270 153798 586302 154034
rect 586538 153798 586622 154034
rect 586858 153798 586890 154034
rect 586270 118354 586890 153798
rect 586270 118118 586302 118354
rect 586538 118118 586622 118354
rect 586858 118118 586890 118354
rect 586270 118034 586890 118118
rect 586270 117798 586302 118034
rect 586538 117798 586622 118034
rect 586858 117798 586890 118034
rect 586270 82354 586890 117798
rect 586270 82118 586302 82354
rect 586538 82118 586622 82354
rect 586858 82118 586890 82354
rect 586270 82034 586890 82118
rect 586270 81798 586302 82034
rect 586538 81798 586622 82034
rect 586858 81798 586890 82034
rect 586270 46354 586890 81798
rect 586270 46118 586302 46354
rect 586538 46118 586622 46354
rect 586858 46118 586890 46354
rect 586270 46034 586890 46118
rect 586270 45798 586302 46034
rect 586538 45798 586622 46034
rect 586858 45798 586890 46034
rect 586270 10354 586890 45798
rect 586270 10118 586302 10354
rect 586538 10118 586622 10354
rect 586858 10118 586890 10354
rect 586270 10034 586890 10118
rect 586270 9798 586302 10034
rect 586538 9798 586622 10034
rect 586858 9798 586890 10034
rect 582294 -1542 582326 -1306
rect 582562 -1542 582646 -1306
rect 582882 -1542 582914 -1306
rect 582294 -1626 582914 -1542
rect 582294 -1862 582326 -1626
rect 582562 -1862 582646 -1626
rect 582882 -1862 582914 -1626
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 582294 -7654 582914 -1862
rect 586270 -1306 586890 9798
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 -2266 587850 706202
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 -3226 588810 707162
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 -4186 589770 708122
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 -5146 590730 709082
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 -6106 591690 710042
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 -7066 592650 711002
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 582326 705562 582562 705798
rect 582646 705562 582882 705798
rect 582326 705242 582562 705478
rect 582646 705242 582882 705478
rect -2934 694118 -2698 694354
rect -2614 694118 -2378 694354
rect -2934 693798 -2698 694034
rect -2614 693798 -2378 694034
rect -2934 658118 -2698 658354
rect -2614 658118 -2378 658354
rect -2934 657798 -2698 658034
rect -2614 657798 -2378 658034
rect -2934 622118 -2698 622354
rect -2614 622118 -2378 622354
rect -2934 621798 -2698 622034
rect -2614 621798 -2378 622034
rect -2934 586118 -2698 586354
rect -2614 586118 -2378 586354
rect -2934 585798 -2698 586034
rect -2614 585798 -2378 586034
rect -2934 550118 -2698 550354
rect -2614 550118 -2378 550354
rect -2934 549798 -2698 550034
rect -2614 549798 -2378 550034
rect -2934 514118 -2698 514354
rect -2614 514118 -2378 514354
rect -2934 513798 -2698 514034
rect -2614 513798 -2378 514034
rect -2934 478118 -2698 478354
rect -2614 478118 -2378 478354
rect -2934 477798 -2698 478034
rect -2614 477798 -2378 478034
rect -2934 442118 -2698 442354
rect -2614 442118 -2378 442354
rect -2934 441798 -2698 442034
rect -2614 441798 -2378 442034
rect -2934 406118 -2698 406354
rect -2614 406118 -2378 406354
rect -2934 405798 -2698 406034
rect -2614 405798 -2378 406034
rect -2934 370118 -2698 370354
rect -2614 370118 -2378 370354
rect -2934 369798 -2698 370034
rect -2614 369798 -2378 370034
rect -2934 334118 -2698 334354
rect -2614 334118 -2378 334354
rect -2934 333798 -2698 334034
rect -2614 333798 -2378 334034
rect -2934 298118 -2698 298354
rect -2614 298118 -2378 298354
rect -2934 297798 -2698 298034
rect -2614 297798 -2378 298034
rect -2934 262118 -2698 262354
rect -2614 262118 -2378 262354
rect -2934 261798 -2698 262034
rect -2614 261798 -2378 262034
rect -2934 226118 -2698 226354
rect -2614 226118 -2378 226354
rect -2934 225798 -2698 226034
rect -2614 225798 -2378 226034
rect -2934 190118 -2698 190354
rect -2614 190118 -2378 190354
rect -2934 189798 -2698 190034
rect -2614 189798 -2378 190034
rect -2934 154118 -2698 154354
rect -2614 154118 -2378 154354
rect -2934 153798 -2698 154034
rect -2614 153798 -2378 154034
rect -2934 118118 -2698 118354
rect -2614 118118 -2378 118354
rect -2934 117798 -2698 118034
rect -2614 117798 -2378 118034
rect -2934 82118 -2698 82354
rect -2614 82118 -2378 82354
rect -2934 81798 -2698 82034
rect -2614 81798 -2378 82034
rect -2934 46118 -2698 46354
rect -2614 46118 -2378 46354
rect -2934 45798 -2698 46034
rect -2614 45798 -2378 46034
rect -2934 10118 -2698 10354
rect -2614 10118 -2378 10354
rect -2934 9798 -2698 10034
rect -2614 9798 -2378 10034
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 23826 694118 24062 694354
rect 24146 694118 24382 694354
rect 23826 693798 24062 694034
rect 24146 693798 24382 694034
rect 59826 694118 60062 694354
rect 60146 694118 60382 694354
rect 59826 693798 60062 694034
rect 60146 693798 60382 694034
rect 95826 694118 96062 694354
rect 96146 694118 96382 694354
rect 95826 693798 96062 694034
rect 96146 693798 96382 694034
rect 131826 694118 132062 694354
rect 132146 694118 132382 694354
rect 131826 693798 132062 694034
rect 132146 693798 132382 694034
rect 167826 694118 168062 694354
rect 168146 694118 168382 694354
rect 167826 693798 168062 694034
rect 168146 693798 168382 694034
rect 203826 694118 204062 694354
rect 204146 694118 204382 694354
rect 203826 693798 204062 694034
rect 204146 693798 204382 694034
rect 239826 694118 240062 694354
rect 240146 694118 240382 694354
rect 239826 693798 240062 694034
rect 240146 693798 240382 694034
rect 275826 694118 276062 694354
rect 276146 694118 276382 694354
rect 275826 693798 276062 694034
rect 276146 693798 276382 694034
rect 311826 694118 312062 694354
rect 312146 694118 312382 694354
rect 311826 693798 312062 694034
rect 312146 693798 312382 694034
rect 347826 694118 348062 694354
rect 348146 694118 348382 694354
rect 347826 693798 348062 694034
rect 348146 693798 348382 694034
rect 383826 694118 384062 694354
rect 384146 694118 384382 694354
rect 383826 693798 384062 694034
rect 384146 693798 384382 694034
rect 419826 694118 420062 694354
rect 420146 694118 420382 694354
rect 419826 693798 420062 694034
rect 420146 693798 420382 694034
rect 455826 694118 456062 694354
rect 456146 694118 456382 694354
rect 455826 693798 456062 694034
rect 456146 693798 456382 694034
rect 491826 694118 492062 694354
rect 492146 694118 492382 694354
rect 491826 693798 492062 694034
rect 492146 693798 492382 694034
rect 527826 694118 528062 694354
rect 528146 694118 528382 694354
rect 527826 693798 528062 694034
rect 528146 693798 528382 694034
rect 563826 694118 564062 694354
rect 564146 694118 564382 694354
rect 563826 693798 564062 694034
rect 564146 693798 564382 694034
rect 582326 694118 582562 694354
rect 582646 694118 582882 694354
rect 582326 693798 582562 694034
rect 582646 693798 582882 694034
rect -1974 689618 -1738 689854
rect -1654 689618 -1418 689854
rect -1974 689298 -1738 689534
rect -1654 689298 -1418 689534
rect 5826 689618 6062 689854
rect 6146 689618 6382 689854
rect 5826 689298 6062 689534
rect 6146 689298 6382 689534
rect 41826 689618 42062 689854
rect 42146 689618 42382 689854
rect 41826 689298 42062 689534
rect 42146 689298 42382 689534
rect 77826 689618 78062 689854
rect 78146 689618 78382 689854
rect 77826 689298 78062 689534
rect 78146 689298 78382 689534
rect 113826 689618 114062 689854
rect 114146 689618 114382 689854
rect 113826 689298 114062 689534
rect 114146 689298 114382 689534
rect 149826 689618 150062 689854
rect 150146 689618 150382 689854
rect 149826 689298 150062 689534
rect 150146 689298 150382 689534
rect 185826 689618 186062 689854
rect 186146 689618 186382 689854
rect 185826 689298 186062 689534
rect 186146 689298 186382 689534
rect 221826 689618 222062 689854
rect 222146 689618 222382 689854
rect 221826 689298 222062 689534
rect 222146 689298 222382 689534
rect 257826 689618 258062 689854
rect 258146 689618 258382 689854
rect 257826 689298 258062 689534
rect 258146 689298 258382 689534
rect 293826 689618 294062 689854
rect 294146 689618 294382 689854
rect 293826 689298 294062 689534
rect 294146 689298 294382 689534
rect 329826 689618 330062 689854
rect 330146 689618 330382 689854
rect 329826 689298 330062 689534
rect 330146 689298 330382 689534
rect 365826 689618 366062 689854
rect 366146 689618 366382 689854
rect 365826 689298 366062 689534
rect 366146 689298 366382 689534
rect 401826 689618 402062 689854
rect 402146 689618 402382 689854
rect 401826 689298 402062 689534
rect 402146 689298 402382 689534
rect 437826 689618 438062 689854
rect 438146 689618 438382 689854
rect 437826 689298 438062 689534
rect 438146 689298 438382 689534
rect 473826 689618 474062 689854
rect 474146 689618 474382 689854
rect 473826 689298 474062 689534
rect 474146 689298 474382 689534
rect 509826 689618 510062 689854
rect 510146 689618 510382 689854
rect 509826 689298 510062 689534
rect 510146 689298 510382 689534
rect 545826 689618 546062 689854
rect 546146 689618 546382 689854
rect 545826 689298 546062 689534
rect 546146 689298 546382 689534
rect 13198 658118 13434 658354
rect 13518 658118 13754 658354
rect 13198 657798 13434 658034
rect 13518 657798 13754 658034
rect 167826 658118 168062 658354
rect 168146 658118 168382 658354
rect 167826 657798 168062 658034
rect 168146 657798 168382 658034
rect 291590 658118 291826 658354
rect 291910 658118 292146 658354
rect 291590 657798 291826 658034
rect 291910 657798 292146 658034
rect 419826 658118 420062 658354
rect 420146 658118 420382 658354
rect 419826 657798 420062 658034
rect 420146 657798 420382 658034
rect 563826 658118 564062 658354
rect 564146 658118 564382 658354
rect 563826 657798 564062 658034
rect 564146 657798 564382 658034
rect 582326 658118 582562 658354
rect 582646 658118 582882 658354
rect 582326 657798 582562 658034
rect 582646 657798 582882 658034
rect -1974 653618 -1738 653854
rect -1654 653618 -1418 653854
rect -1974 653298 -1738 653534
rect -1654 653298 -1418 653534
rect 5826 653618 6062 653854
rect 6146 653618 6382 653854
rect 5826 653298 6062 653534
rect 6146 653298 6382 653534
rect 173094 653618 173330 653854
rect 173414 653618 173650 653854
rect 173094 653298 173330 653534
rect 173414 653298 173650 653534
rect 293826 653618 294062 653854
rect 294146 653618 294382 653854
rect 293826 653298 294062 653534
rect 294146 653298 294382 653534
rect 401826 653618 402062 653854
rect 402146 653618 402382 653854
rect 401826 653298 402062 653534
rect 402146 653298 402382 653534
rect 570350 653618 570586 653854
rect 570670 653618 570906 653854
rect 570350 653298 570586 653534
rect 570670 653298 570906 653534
rect 13198 622118 13434 622354
rect 13518 622118 13754 622354
rect 13198 621798 13434 622034
rect 13518 621798 13754 622034
rect 167826 622118 168062 622354
rect 168146 622118 168382 622354
rect 167826 621798 168062 622034
rect 168146 621798 168382 622034
rect 291590 622118 291826 622354
rect 291910 622118 292146 622354
rect 291590 621798 291826 622034
rect 291910 621798 292146 622034
rect 419826 622118 420062 622354
rect 420146 622118 420382 622354
rect 419826 621798 420062 622034
rect 420146 621798 420382 622034
rect 563826 622118 564062 622354
rect 564146 622118 564382 622354
rect 563826 621798 564062 622034
rect 564146 621798 564382 622034
rect 582326 622118 582562 622354
rect 582646 622118 582882 622354
rect 582326 621798 582562 622034
rect 582646 621798 582882 622034
rect -1974 617618 -1738 617854
rect -1654 617618 -1418 617854
rect -1974 617298 -1738 617534
rect -1654 617298 -1418 617534
rect 5826 617618 6062 617854
rect 6146 617618 6382 617854
rect 5826 617298 6062 617534
rect 6146 617298 6382 617534
rect 173094 617618 173330 617854
rect 173414 617618 173650 617854
rect 173094 617298 173330 617534
rect 173414 617298 173650 617534
rect 293826 617618 294062 617854
rect 294146 617618 294382 617854
rect 293826 617298 294062 617534
rect 294146 617298 294382 617534
rect 401826 617618 402062 617854
rect 402146 617618 402382 617854
rect 401826 617298 402062 617534
rect 402146 617298 402382 617534
rect 570350 617618 570586 617854
rect 570670 617618 570906 617854
rect 570350 617298 570586 617534
rect 570670 617298 570906 617534
rect 23826 586118 24062 586354
rect 24146 586118 24382 586354
rect 23826 585798 24062 586034
rect 24146 585798 24382 586034
rect 59826 586118 60062 586354
rect 60146 586118 60382 586354
rect 59826 585798 60062 586034
rect 60146 585798 60382 586034
rect 95826 586118 96062 586354
rect 96146 586118 96382 586354
rect 95826 585798 96062 586034
rect 96146 585798 96382 586034
rect 131826 586118 132062 586354
rect 132146 586118 132382 586354
rect 131826 585798 132062 586034
rect 132146 585798 132382 586034
rect 167826 586118 168062 586354
rect 168146 586118 168382 586354
rect 167826 585798 168062 586034
rect 168146 585798 168382 586034
rect 203826 586118 204062 586354
rect 204146 586118 204382 586354
rect 203826 585798 204062 586034
rect 204146 585798 204382 586034
rect 239826 586118 240062 586354
rect 240146 586118 240382 586354
rect 239826 585798 240062 586034
rect 240146 585798 240382 586034
rect 275826 586118 276062 586354
rect 276146 586118 276382 586354
rect 275826 585798 276062 586034
rect 276146 585798 276382 586034
rect 311826 586118 312062 586354
rect 312146 586118 312382 586354
rect 311826 585798 312062 586034
rect 312146 585798 312382 586034
rect 347826 586118 348062 586354
rect 348146 586118 348382 586354
rect 347826 585798 348062 586034
rect 348146 585798 348382 586034
rect 383826 586118 384062 586354
rect 384146 586118 384382 586354
rect 383826 585798 384062 586034
rect 384146 585798 384382 586034
rect 419826 586118 420062 586354
rect 420146 586118 420382 586354
rect 419826 585798 420062 586034
rect 420146 585798 420382 586034
rect 455826 586118 456062 586354
rect 456146 586118 456382 586354
rect 455826 585798 456062 586034
rect 456146 585798 456382 586034
rect 491826 586118 492062 586354
rect 492146 586118 492382 586354
rect 491826 585798 492062 586034
rect 492146 585798 492382 586034
rect 527826 586118 528062 586354
rect 528146 586118 528382 586354
rect 527826 585798 528062 586034
rect 528146 585798 528382 586034
rect 563826 586118 564062 586354
rect 564146 586118 564382 586354
rect 563826 585798 564062 586034
rect 564146 585798 564382 586034
rect 582326 586118 582562 586354
rect 582646 586118 582882 586354
rect 582326 585798 582562 586034
rect 582646 585798 582882 586034
rect -1974 581618 -1738 581854
rect -1654 581618 -1418 581854
rect -1974 581298 -1738 581534
rect -1654 581298 -1418 581534
rect 5826 581618 6062 581854
rect 6146 581618 6382 581854
rect 5826 581298 6062 581534
rect 6146 581298 6382 581534
rect 41826 581618 42062 581854
rect 42146 581618 42382 581854
rect 41826 581298 42062 581534
rect 42146 581298 42382 581534
rect 77826 581618 78062 581854
rect 78146 581618 78382 581854
rect 77826 581298 78062 581534
rect 78146 581298 78382 581534
rect 113826 581618 114062 581854
rect 114146 581618 114382 581854
rect 113826 581298 114062 581534
rect 114146 581298 114382 581534
rect 149826 581618 150062 581854
rect 150146 581618 150382 581854
rect 149826 581298 150062 581534
rect 150146 581298 150382 581534
rect 185826 581618 186062 581854
rect 186146 581618 186382 581854
rect 185826 581298 186062 581534
rect 186146 581298 186382 581534
rect 221826 581618 222062 581854
rect 222146 581618 222382 581854
rect 221826 581298 222062 581534
rect 222146 581298 222382 581534
rect 257826 581618 258062 581854
rect 258146 581618 258382 581854
rect 257826 581298 258062 581534
rect 258146 581298 258382 581534
rect 293826 581618 294062 581854
rect 294146 581618 294382 581854
rect 293826 581298 294062 581534
rect 294146 581298 294382 581534
rect 329826 581618 330062 581854
rect 330146 581618 330382 581854
rect 329826 581298 330062 581534
rect 330146 581298 330382 581534
rect 365826 581618 366062 581854
rect 366146 581618 366382 581854
rect 365826 581298 366062 581534
rect 366146 581298 366382 581534
rect 401826 581618 402062 581854
rect 402146 581618 402382 581854
rect 401826 581298 402062 581534
rect 402146 581298 402382 581534
rect 437826 581618 438062 581854
rect 438146 581618 438382 581854
rect 437826 581298 438062 581534
rect 438146 581298 438382 581534
rect 473826 581618 474062 581854
rect 474146 581618 474382 581854
rect 473826 581298 474062 581534
rect 474146 581298 474382 581534
rect 509826 581618 510062 581854
rect 510146 581618 510382 581854
rect 509826 581298 510062 581534
rect 510146 581298 510382 581534
rect 545826 581618 546062 581854
rect 546146 581618 546382 581854
rect 545826 581298 546062 581534
rect 546146 581298 546382 581534
rect 13198 550118 13434 550354
rect 13518 550118 13754 550354
rect 13198 549798 13434 550034
rect 13518 549798 13754 550034
rect 167826 550118 168062 550354
rect 168146 550118 168382 550354
rect 167826 549798 168062 550034
rect 168146 549798 168382 550034
rect 203826 550118 204062 550354
rect 204146 550118 204382 550354
rect 203826 549798 204062 550034
rect 204146 549798 204382 550034
rect 239826 550118 240062 550354
rect 240146 550118 240382 550354
rect 239826 549798 240062 550034
rect 240146 549798 240382 550034
rect 275826 550118 276062 550354
rect 276146 550118 276382 550354
rect 275826 549798 276062 550034
rect 276146 549798 276382 550034
rect 311826 550118 312062 550354
rect 312146 550118 312382 550354
rect 311826 549798 312062 550034
rect 312146 549798 312382 550034
rect 347826 550118 348062 550354
rect 348146 550118 348382 550354
rect 347826 549798 348062 550034
rect 348146 549798 348382 550034
rect 383826 550118 384062 550354
rect 384146 550118 384382 550354
rect 383826 549798 384062 550034
rect 384146 549798 384382 550034
rect 419826 550118 420062 550354
rect 420146 550118 420382 550354
rect 419826 549798 420062 550034
rect 420146 549798 420382 550034
rect 563826 550118 564062 550354
rect 564146 550118 564382 550354
rect 563826 549798 564062 550034
rect 564146 549798 564382 550034
rect 582326 550118 582562 550354
rect 582646 550118 582882 550354
rect 582326 549798 582562 550034
rect 582646 549798 582882 550034
rect -1974 545618 -1738 545854
rect -1654 545618 -1418 545854
rect -1974 545298 -1738 545534
rect -1654 545298 -1418 545534
rect 5826 545618 6062 545854
rect 6146 545618 6382 545854
rect 5826 545298 6062 545534
rect 6146 545298 6382 545534
rect 185826 545618 186062 545854
rect 186146 545618 186382 545854
rect 185826 545298 186062 545534
rect 186146 545298 186382 545534
rect 221826 545618 222062 545854
rect 222146 545618 222382 545854
rect 221826 545298 222062 545534
rect 222146 545298 222382 545534
rect 257826 545618 258062 545854
rect 258146 545618 258382 545854
rect 257826 545298 258062 545534
rect 258146 545298 258382 545534
rect 293826 545618 294062 545854
rect 294146 545618 294382 545854
rect 293826 545298 294062 545534
rect 294146 545298 294382 545534
rect 329826 545618 330062 545854
rect 330146 545618 330382 545854
rect 329826 545298 330062 545534
rect 330146 545298 330382 545534
rect 365826 545618 366062 545854
rect 366146 545618 366382 545854
rect 365826 545298 366062 545534
rect 366146 545298 366382 545534
rect 401826 545618 402062 545854
rect 402146 545618 402382 545854
rect 401826 545298 402062 545534
rect 402146 545298 402382 545534
rect 570350 545618 570586 545854
rect 570670 545618 570906 545854
rect 570350 545298 570586 545534
rect 570670 545298 570906 545534
rect 13198 514118 13434 514354
rect 13518 514118 13754 514354
rect 13198 513798 13434 514034
rect 13518 513798 13754 514034
rect 167826 514118 168062 514354
rect 168146 514118 168382 514354
rect 167826 513798 168062 514034
rect 168146 513798 168382 514034
rect 203826 514118 204062 514354
rect 204146 514118 204382 514354
rect 203826 513798 204062 514034
rect 204146 513798 204382 514034
rect 239826 514118 240062 514354
rect 240146 514118 240382 514354
rect 239826 513798 240062 514034
rect 240146 513798 240382 514034
rect 275826 514118 276062 514354
rect 276146 514118 276382 514354
rect 275826 513798 276062 514034
rect 276146 513798 276382 514034
rect 311826 514118 312062 514354
rect 312146 514118 312382 514354
rect 311826 513798 312062 514034
rect 312146 513798 312382 514034
rect 347826 514118 348062 514354
rect 348146 514118 348382 514354
rect 347826 513798 348062 514034
rect 348146 513798 348382 514034
rect 383826 514118 384062 514354
rect 384146 514118 384382 514354
rect 383826 513798 384062 514034
rect 384146 513798 384382 514034
rect 419826 514118 420062 514354
rect 420146 514118 420382 514354
rect 419826 513798 420062 514034
rect 420146 513798 420382 514034
rect 563826 514118 564062 514354
rect 564146 514118 564382 514354
rect 563826 513798 564062 514034
rect 564146 513798 564382 514034
rect 582326 514118 582562 514354
rect 582646 514118 582882 514354
rect 582326 513798 582562 514034
rect 582646 513798 582882 514034
rect -1974 509618 -1738 509854
rect -1654 509618 -1418 509854
rect -1974 509298 -1738 509534
rect -1654 509298 -1418 509534
rect 5826 509618 6062 509854
rect 6146 509618 6382 509854
rect 5826 509298 6062 509534
rect 6146 509298 6382 509534
rect 185826 509618 186062 509854
rect 186146 509618 186382 509854
rect 185826 509298 186062 509534
rect 186146 509298 186382 509534
rect 221826 509618 222062 509854
rect 222146 509618 222382 509854
rect 221826 509298 222062 509534
rect 222146 509298 222382 509534
rect 257826 509618 258062 509854
rect 258146 509618 258382 509854
rect 257826 509298 258062 509534
rect 258146 509298 258382 509534
rect 293826 509618 294062 509854
rect 294146 509618 294382 509854
rect 293826 509298 294062 509534
rect 294146 509298 294382 509534
rect 329826 509618 330062 509854
rect 330146 509618 330382 509854
rect 329826 509298 330062 509534
rect 330146 509298 330382 509534
rect 365826 509618 366062 509854
rect 366146 509618 366382 509854
rect 365826 509298 366062 509534
rect 366146 509298 366382 509534
rect 401826 509618 402062 509854
rect 402146 509618 402382 509854
rect 401826 509298 402062 509534
rect 402146 509298 402382 509534
rect 570350 509618 570586 509854
rect 570670 509618 570906 509854
rect 570350 509298 570586 509534
rect 570670 509298 570906 509534
rect 23826 478118 24062 478354
rect 24146 478118 24382 478354
rect 23826 477798 24062 478034
rect 24146 477798 24382 478034
rect 59826 478118 60062 478354
rect 60146 478118 60382 478354
rect 59826 477798 60062 478034
rect 60146 477798 60382 478034
rect 95826 478118 96062 478354
rect 96146 478118 96382 478354
rect 95826 477798 96062 478034
rect 96146 477798 96382 478034
rect 131826 478118 132062 478354
rect 132146 478118 132382 478354
rect 131826 477798 132062 478034
rect 132146 477798 132382 478034
rect 167826 478118 168062 478354
rect 168146 478118 168382 478354
rect 167826 477798 168062 478034
rect 168146 477798 168382 478034
rect 203826 478118 204062 478354
rect 204146 478118 204382 478354
rect 203826 477798 204062 478034
rect 204146 477798 204382 478034
rect 239826 478118 240062 478354
rect 240146 478118 240382 478354
rect 239826 477798 240062 478034
rect 240146 477798 240382 478034
rect 275826 478118 276062 478354
rect 276146 478118 276382 478354
rect 275826 477798 276062 478034
rect 276146 477798 276382 478034
rect 311826 478118 312062 478354
rect 312146 478118 312382 478354
rect 311826 477798 312062 478034
rect 312146 477798 312382 478034
rect 347826 478118 348062 478354
rect 348146 478118 348382 478354
rect 347826 477798 348062 478034
rect 348146 477798 348382 478034
rect 383826 478118 384062 478354
rect 384146 478118 384382 478354
rect 383826 477798 384062 478034
rect 384146 477798 384382 478034
rect 419826 478118 420062 478354
rect 420146 478118 420382 478354
rect 419826 477798 420062 478034
rect 420146 477798 420382 478034
rect 455826 478118 456062 478354
rect 456146 478118 456382 478354
rect 455826 477798 456062 478034
rect 456146 477798 456382 478034
rect 491826 478118 492062 478354
rect 492146 478118 492382 478354
rect 491826 477798 492062 478034
rect 492146 477798 492382 478034
rect 527826 478118 528062 478354
rect 528146 478118 528382 478354
rect 527826 477798 528062 478034
rect 528146 477798 528382 478034
rect 563826 478118 564062 478354
rect 564146 478118 564382 478354
rect 563826 477798 564062 478034
rect 564146 477798 564382 478034
rect 582326 478118 582562 478354
rect 582646 478118 582882 478354
rect 582326 477798 582562 478034
rect 582646 477798 582882 478034
rect -1974 473618 -1738 473854
rect -1654 473618 -1418 473854
rect -1974 473298 -1738 473534
rect -1654 473298 -1418 473534
rect 5826 473618 6062 473854
rect 6146 473618 6382 473854
rect 5826 473298 6062 473534
rect 6146 473298 6382 473534
rect 41826 473618 42062 473854
rect 42146 473618 42382 473854
rect 41826 473298 42062 473534
rect 42146 473298 42382 473534
rect 77826 473618 78062 473854
rect 78146 473618 78382 473854
rect 77826 473298 78062 473534
rect 78146 473298 78382 473534
rect 113826 473618 114062 473854
rect 114146 473618 114382 473854
rect 113826 473298 114062 473534
rect 114146 473298 114382 473534
rect 149826 473618 150062 473854
rect 150146 473618 150382 473854
rect 149826 473298 150062 473534
rect 150146 473298 150382 473534
rect 185826 473618 186062 473854
rect 186146 473618 186382 473854
rect 185826 473298 186062 473534
rect 186146 473298 186382 473534
rect 221826 473618 222062 473854
rect 222146 473618 222382 473854
rect 221826 473298 222062 473534
rect 222146 473298 222382 473534
rect 257826 473618 258062 473854
rect 258146 473618 258382 473854
rect 257826 473298 258062 473534
rect 258146 473298 258382 473534
rect 293826 473618 294062 473854
rect 294146 473618 294382 473854
rect 293826 473298 294062 473534
rect 294146 473298 294382 473534
rect 329826 473618 330062 473854
rect 330146 473618 330382 473854
rect 329826 473298 330062 473534
rect 330146 473298 330382 473534
rect 365826 473618 366062 473854
rect 366146 473618 366382 473854
rect 365826 473298 366062 473534
rect 366146 473298 366382 473534
rect 401826 473618 402062 473854
rect 402146 473618 402382 473854
rect 401826 473298 402062 473534
rect 402146 473298 402382 473534
rect 437826 473618 438062 473854
rect 438146 473618 438382 473854
rect 437826 473298 438062 473534
rect 438146 473298 438382 473534
rect 473826 473618 474062 473854
rect 474146 473618 474382 473854
rect 473826 473298 474062 473534
rect 474146 473298 474382 473534
rect 509826 473618 510062 473854
rect 510146 473618 510382 473854
rect 509826 473298 510062 473534
rect 510146 473298 510382 473534
rect 545826 473618 546062 473854
rect 546146 473618 546382 473854
rect 545826 473298 546062 473534
rect 546146 473298 546382 473534
rect 13198 442118 13434 442354
rect 13518 442118 13754 442354
rect 13198 441798 13434 442034
rect 13518 441798 13754 442034
rect 167826 442118 168062 442354
rect 168146 442118 168382 442354
rect 167826 441798 168062 442034
rect 168146 441798 168382 442034
rect 203826 442118 204062 442354
rect 204146 442118 204382 442354
rect 203826 441798 204062 442034
rect 204146 441798 204382 442034
rect 239826 442118 240062 442354
rect 240146 442118 240382 442354
rect 239826 441798 240062 442034
rect 240146 441798 240382 442034
rect 275826 442118 276062 442354
rect 276146 442118 276382 442354
rect 275826 441798 276062 442034
rect 276146 441798 276382 442034
rect 311826 442118 312062 442354
rect 312146 442118 312382 442354
rect 311826 441798 312062 442034
rect 312146 441798 312382 442034
rect 347826 442118 348062 442354
rect 348146 442118 348382 442354
rect 347826 441798 348062 442034
rect 348146 441798 348382 442034
rect 383826 442118 384062 442354
rect 384146 442118 384382 442354
rect 383826 441798 384062 442034
rect 384146 441798 384382 442034
rect 419826 442118 420062 442354
rect 420146 442118 420382 442354
rect 419826 441798 420062 442034
rect 420146 441798 420382 442034
rect 563826 442118 564062 442354
rect 564146 442118 564382 442354
rect 563826 441798 564062 442034
rect 564146 441798 564382 442034
rect 582326 442118 582562 442354
rect 582646 442118 582882 442354
rect 582326 441798 582562 442034
rect 582646 441798 582882 442034
rect -1974 437618 -1738 437854
rect -1654 437618 -1418 437854
rect -1974 437298 -1738 437534
rect -1654 437298 -1418 437534
rect 5826 437618 6062 437854
rect 6146 437618 6382 437854
rect 5826 437298 6062 437534
rect 6146 437298 6382 437534
rect 185826 437618 186062 437854
rect 186146 437618 186382 437854
rect 185826 437298 186062 437534
rect 186146 437298 186382 437534
rect 221826 437618 222062 437854
rect 222146 437618 222382 437854
rect 221826 437298 222062 437534
rect 222146 437298 222382 437534
rect 257826 437618 258062 437854
rect 258146 437618 258382 437854
rect 257826 437298 258062 437534
rect 258146 437298 258382 437534
rect 293826 437618 294062 437854
rect 294146 437618 294382 437854
rect 293826 437298 294062 437534
rect 294146 437298 294382 437534
rect 329826 437618 330062 437854
rect 330146 437618 330382 437854
rect 329826 437298 330062 437534
rect 330146 437298 330382 437534
rect 365826 437618 366062 437854
rect 366146 437618 366382 437854
rect 365826 437298 366062 437534
rect 366146 437298 366382 437534
rect 401826 437618 402062 437854
rect 402146 437618 402382 437854
rect 401826 437298 402062 437534
rect 402146 437298 402382 437534
rect 570350 437618 570586 437854
rect 570670 437618 570906 437854
rect 570350 437298 570586 437534
rect 570670 437298 570906 437534
rect 13198 406118 13434 406354
rect 13518 406118 13754 406354
rect 13198 405798 13434 406034
rect 13518 405798 13754 406034
rect 167826 406118 168062 406354
rect 168146 406118 168382 406354
rect 167826 405798 168062 406034
rect 168146 405798 168382 406034
rect 203826 406118 204062 406354
rect 204146 406118 204382 406354
rect 203826 405798 204062 406034
rect 204146 405798 204382 406034
rect 239826 406118 240062 406354
rect 240146 406118 240382 406354
rect 239826 405798 240062 406034
rect 240146 405798 240382 406034
rect 275826 406118 276062 406354
rect 276146 406118 276382 406354
rect 275826 405798 276062 406034
rect 276146 405798 276382 406034
rect 311826 406118 312062 406354
rect 312146 406118 312382 406354
rect 311826 405798 312062 406034
rect 312146 405798 312382 406034
rect 347826 406118 348062 406354
rect 348146 406118 348382 406354
rect 347826 405798 348062 406034
rect 348146 405798 348382 406034
rect 383826 406118 384062 406354
rect 384146 406118 384382 406354
rect 383826 405798 384062 406034
rect 384146 405798 384382 406034
rect 419826 406118 420062 406354
rect 420146 406118 420382 406354
rect 419826 405798 420062 406034
rect 420146 405798 420382 406034
rect 563826 406118 564062 406354
rect 564146 406118 564382 406354
rect 563826 405798 564062 406034
rect 564146 405798 564382 406034
rect 582326 406118 582562 406354
rect 582646 406118 582882 406354
rect 582326 405798 582562 406034
rect 582646 405798 582882 406034
rect -1974 401618 -1738 401854
rect -1654 401618 -1418 401854
rect -1974 401298 -1738 401534
rect -1654 401298 -1418 401534
rect 5826 401618 6062 401854
rect 6146 401618 6382 401854
rect 5826 401298 6062 401534
rect 6146 401298 6382 401534
rect 185826 401618 186062 401854
rect 186146 401618 186382 401854
rect 185826 401298 186062 401534
rect 186146 401298 186382 401534
rect 221826 401618 222062 401854
rect 222146 401618 222382 401854
rect 221826 401298 222062 401534
rect 222146 401298 222382 401534
rect 257826 401618 258062 401854
rect 258146 401618 258382 401854
rect 257826 401298 258062 401534
rect 258146 401298 258382 401534
rect 293826 401618 294062 401854
rect 294146 401618 294382 401854
rect 293826 401298 294062 401534
rect 294146 401298 294382 401534
rect 329826 401618 330062 401854
rect 330146 401618 330382 401854
rect 329826 401298 330062 401534
rect 330146 401298 330382 401534
rect 365826 401618 366062 401854
rect 366146 401618 366382 401854
rect 365826 401298 366062 401534
rect 366146 401298 366382 401534
rect 401826 401618 402062 401854
rect 402146 401618 402382 401854
rect 401826 401298 402062 401534
rect 402146 401298 402382 401534
rect 570350 401618 570586 401854
rect 570670 401618 570906 401854
rect 570350 401298 570586 401534
rect 570670 401298 570906 401534
rect 13198 370118 13434 370354
rect 13518 370118 13754 370354
rect 13198 369798 13434 370034
rect 13518 369798 13754 370034
rect 167826 370118 168062 370354
rect 168146 370118 168382 370354
rect 167826 369798 168062 370034
rect 168146 369798 168382 370034
rect 203826 370118 204062 370354
rect 204146 370118 204382 370354
rect 203826 369798 204062 370034
rect 204146 369798 204382 370034
rect 239826 370118 240062 370354
rect 240146 370118 240382 370354
rect 239826 369798 240062 370034
rect 240146 369798 240382 370034
rect 275826 370118 276062 370354
rect 276146 370118 276382 370354
rect 275826 369798 276062 370034
rect 276146 369798 276382 370034
rect 311826 370118 312062 370354
rect 312146 370118 312382 370354
rect 311826 369798 312062 370034
rect 312146 369798 312382 370034
rect 347826 370118 348062 370354
rect 348146 370118 348382 370354
rect 347826 369798 348062 370034
rect 348146 369798 348382 370034
rect 383826 370118 384062 370354
rect 384146 370118 384382 370354
rect 383826 369798 384062 370034
rect 384146 369798 384382 370034
rect 419826 370118 420062 370354
rect 420146 370118 420382 370354
rect 419826 369798 420062 370034
rect 420146 369798 420382 370034
rect 563826 370118 564062 370354
rect 564146 370118 564382 370354
rect 563826 369798 564062 370034
rect 564146 369798 564382 370034
rect 582326 370118 582562 370354
rect 582646 370118 582882 370354
rect 582326 369798 582562 370034
rect 582646 369798 582882 370034
rect -1974 365618 -1738 365854
rect -1654 365618 -1418 365854
rect -1974 365298 -1738 365534
rect -1654 365298 -1418 365534
rect 5826 365618 6062 365854
rect 6146 365618 6382 365854
rect 5826 365298 6062 365534
rect 6146 365298 6382 365534
rect 41826 365618 42062 365854
rect 42146 365618 42382 365854
rect 41826 365298 42062 365534
rect 42146 365298 42382 365534
rect 77826 365618 78062 365854
rect 78146 365618 78382 365854
rect 77826 365298 78062 365534
rect 78146 365298 78382 365534
rect 113826 365618 114062 365854
rect 114146 365618 114382 365854
rect 113826 365298 114062 365534
rect 114146 365298 114382 365534
rect 149826 365618 150062 365854
rect 150146 365618 150382 365854
rect 149826 365298 150062 365534
rect 150146 365298 150382 365534
rect 185826 365618 186062 365854
rect 186146 365618 186382 365854
rect 185826 365298 186062 365534
rect 186146 365298 186382 365534
rect 221826 365618 222062 365854
rect 222146 365618 222382 365854
rect 221826 365298 222062 365534
rect 222146 365298 222382 365534
rect 257826 365618 258062 365854
rect 258146 365618 258382 365854
rect 257826 365298 258062 365534
rect 258146 365298 258382 365534
rect 293826 365618 294062 365854
rect 294146 365618 294382 365854
rect 293826 365298 294062 365534
rect 294146 365298 294382 365534
rect 329826 365618 330062 365854
rect 330146 365618 330382 365854
rect 329826 365298 330062 365534
rect 330146 365298 330382 365534
rect 365826 365618 366062 365854
rect 366146 365618 366382 365854
rect 365826 365298 366062 365534
rect 366146 365298 366382 365534
rect 401826 365618 402062 365854
rect 402146 365618 402382 365854
rect 401826 365298 402062 365534
rect 402146 365298 402382 365534
rect 437826 365618 438062 365854
rect 438146 365618 438382 365854
rect 437826 365298 438062 365534
rect 438146 365298 438382 365534
rect 473826 365618 474062 365854
rect 474146 365618 474382 365854
rect 473826 365298 474062 365534
rect 474146 365298 474382 365534
rect 509826 365618 510062 365854
rect 510146 365618 510382 365854
rect 509826 365298 510062 365534
rect 510146 365298 510382 365534
rect 545826 365618 546062 365854
rect 546146 365618 546382 365854
rect 545826 365298 546062 365534
rect 546146 365298 546382 365534
rect 13198 334118 13434 334354
rect 13518 334118 13754 334354
rect 13198 333798 13434 334034
rect 13518 333798 13754 334034
rect 167826 334118 168062 334354
rect 168146 334118 168382 334354
rect 167826 333798 168062 334034
rect 168146 333798 168382 334034
rect 203826 334118 204062 334354
rect 204146 334118 204382 334354
rect 203826 333798 204062 334034
rect 204146 333798 204382 334034
rect 239826 334118 240062 334354
rect 240146 334118 240382 334354
rect 239826 333798 240062 334034
rect 240146 333798 240382 334034
rect 275826 334118 276062 334354
rect 276146 334118 276382 334354
rect 275826 333798 276062 334034
rect 276146 333798 276382 334034
rect 311826 334118 312062 334354
rect 312146 334118 312382 334354
rect 311826 333798 312062 334034
rect 312146 333798 312382 334034
rect 347826 334118 348062 334354
rect 348146 334118 348382 334354
rect 347826 333798 348062 334034
rect 348146 333798 348382 334034
rect 383826 334118 384062 334354
rect 384146 334118 384382 334354
rect 383826 333798 384062 334034
rect 384146 333798 384382 334034
rect 419826 334118 420062 334354
rect 420146 334118 420382 334354
rect 419826 333798 420062 334034
rect 420146 333798 420382 334034
rect 563826 334118 564062 334354
rect 564146 334118 564382 334354
rect 563826 333798 564062 334034
rect 564146 333798 564382 334034
rect 582326 334118 582562 334354
rect 582646 334118 582882 334354
rect 582326 333798 582562 334034
rect 582646 333798 582882 334034
rect -1974 329618 -1738 329854
rect -1654 329618 -1418 329854
rect -1974 329298 -1738 329534
rect -1654 329298 -1418 329534
rect 5826 329618 6062 329854
rect 6146 329618 6382 329854
rect 5826 329298 6062 329534
rect 6146 329298 6382 329534
rect 185826 329618 186062 329854
rect 186146 329618 186382 329854
rect 185826 329298 186062 329534
rect 186146 329298 186382 329534
rect 221826 329618 222062 329854
rect 222146 329618 222382 329854
rect 221826 329298 222062 329534
rect 222146 329298 222382 329534
rect 257826 329618 258062 329854
rect 258146 329618 258382 329854
rect 257826 329298 258062 329534
rect 258146 329298 258382 329534
rect 293826 329618 294062 329854
rect 294146 329618 294382 329854
rect 293826 329298 294062 329534
rect 294146 329298 294382 329534
rect 329826 329618 330062 329854
rect 330146 329618 330382 329854
rect 329826 329298 330062 329534
rect 330146 329298 330382 329534
rect 365826 329618 366062 329854
rect 366146 329618 366382 329854
rect 365826 329298 366062 329534
rect 366146 329298 366382 329534
rect 401826 329618 402062 329854
rect 402146 329618 402382 329854
rect 401826 329298 402062 329534
rect 402146 329298 402382 329534
rect 570350 329618 570586 329854
rect 570670 329618 570906 329854
rect 570350 329298 570586 329534
rect 570670 329298 570906 329534
rect 13198 298118 13434 298354
rect 13518 298118 13754 298354
rect 13198 297798 13434 298034
rect 13518 297798 13754 298034
rect 167826 298118 168062 298354
rect 168146 298118 168382 298354
rect 167826 297798 168062 298034
rect 168146 297798 168382 298034
rect 203826 298118 204062 298354
rect 204146 298118 204382 298354
rect 203826 297798 204062 298034
rect 204146 297798 204382 298034
rect 239826 298118 240062 298354
rect 240146 298118 240382 298354
rect 239826 297798 240062 298034
rect 240146 297798 240382 298034
rect 275826 298118 276062 298354
rect 276146 298118 276382 298354
rect 275826 297798 276062 298034
rect 276146 297798 276382 298034
rect 311826 298118 312062 298354
rect 312146 298118 312382 298354
rect 311826 297798 312062 298034
rect 312146 297798 312382 298034
rect 347826 298118 348062 298354
rect 348146 298118 348382 298354
rect 347826 297798 348062 298034
rect 348146 297798 348382 298034
rect 383826 298118 384062 298354
rect 384146 298118 384382 298354
rect 383826 297798 384062 298034
rect 384146 297798 384382 298034
rect 419826 298118 420062 298354
rect 420146 298118 420382 298354
rect 419826 297798 420062 298034
rect 420146 297798 420382 298034
rect 563826 298118 564062 298354
rect 564146 298118 564382 298354
rect 563826 297798 564062 298034
rect 564146 297798 564382 298034
rect 582326 298118 582562 298354
rect 582646 298118 582882 298354
rect 582326 297798 582562 298034
rect 582646 297798 582882 298034
rect -1974 293618 -1738 293854
rect -1654 293618 -1418 293854
rect -1974 293298 -1738 293534
rect -1654 293298 -1418 293534
rect 5826 293618 6062 293854
rect 6146 293618 6382 293854
rect 5826 293298 6062 293534
rect 6146 293298 6382 293534
rect 185826 293618 186062 293854
rect 186146 293618 186382 293854
rect 185826 293298 186062 293534
rect 186146 293298 186382 293534
rect 221826 293618 222062 293854
rect 222146 293618 222382 293854
rect 221826 293298 222062 293534
rect 222146 293298 222382 293534
rect 257826 293618 258062 293854
rect 258146 293618 258382 293854
rect 257826 293298 258062 293534
rect 258146 293298 258382 293534
rect 293826 293618 294062 293854
rect 294146 293618 294382 293854
rect 293826 293298 294062 293534
rect 294146 293298 294382 293534
rect 329826 293618 330062 293854
rect 330146 293618 330382 293854
rect 329826 293298 330062 293534
rect 330146 293298 330382 293534
rect 365826 293618 366062 293854
rect 366146 293618 366382 293854
rect 365826 293298 366062 293534
rect 366146 293298 366382 293534
rect 401826 293618 402062 293854
rect 402146 293618 402382 293854
rect 401826 293298 402062 293534
rect 402146 293298 402382 293534
rect 570350 293618 570586 293854
rect 570670 293618 570906 293854
rect 570350 293298 570586 293534
rect 570670 293298 570906 293534
rect 13198 262118 13434 262354
rect 13518 262118 13754 262354
rect 13198 261798 13434 262034
rect 13518 261798 13754 262034
rect 167826 262118 168062 262354
rect 168146 262118 168382 262354
rect 167826 261798 168062 262034
rect 168146 261798 168382 262034
rect 203826 262118 204062 262354
rect 204146 262118 204382 262354
rect 203826 261798 204062 262034
rect 204146 261798 204382 262034
rect 239826 262118 240062 262354
rect 240146 262118 240382 262354
rect 239826 261798 240062 262034
rect 240146 261798 240382 262034
rect 275826 262118 276062 262354
rect 276146 262118 276382 262354
rect 275826 261798 276062 262034
rect 276146 261798 276382 262034
rect 311826 262118 312062 262354
rect 312146 262118 312382 262354
rect 311826 261798 312062 262034
rect 312146 261798 312382 262034
rect 347826 262118 348062 262354
rect 348146 262118 348382 262354
rect 347826 261798 348062 262034
rect 348146 261798 348382 262034
rect 383826 262118 384062 262354
rect 384146 262118 384382 262354
rect 383826 261798 384062 262034
rect 384146 261798 384382 262034
rect 419826 262118 420062 262354
rect 420146 262118 420382 262354
rect 419826 261798 420062 262034
rect 420146 261798 420382 262034
rect 563826 262118 564062 262354
rect 564146 262118 564382 262354
rect 563826 261798 564062 262034
rect 564146 261798 564382 262034
rect 582326 262118 582562 262354
rect 582646 262118 582882 262354
rect 582326 261798 582562 262034
rect 582646 261798 582882 262034
rect -1974 257618 -1738 257854
rect -1654 257618 -1418 257854
rect -1974 257298 -1738 257534
rect -1654 257298 -1418 257534
rect 5826 257618 6062 257854
rect 6146 257618 6382 257854
rect 5826 257298 6062 257534
rect 6146 257298 6382 257534
rect 185826 257618 186062 257854
rect 186146 257618 186382 257854
rect 185826 257298 186062 257534
rect 186146 257298 186382 257534
rect 221826 257618 222062 257854
rect 222146 257618 222382 257854
rect 221826 257298 222062 257534
rect 222146 257298 222382 257534
rect 257826 257618 258062 257854
rect 258146 257618 258382 257854
rect 257826 257298 258062 257534
rect 258146 257298 258382 257534
rect 293826 257618 294062 257854
rect 294146 257618 294382 257854
rect 293826 257298 294062 257534
rect 294146 257298 294382 257534
rect 329826 257618 330062 257854
rect 330146 257618 330382 257854
rect 329826 257298 330062 257534
rect 330146 257298 330382 257534
rect 365826 257618 366062 257854
rect 366146 257618 366382 257854
rect 365826 257298 366062 257534
rect 366146 257298 366382 257534
rect 401826 257618 402062 257854
rect 402146 257618 402382 257854
rect 401826 257298 402062 257534
rect 402146 257298 402382 257534
rect 570350 257618 570586 257854
rect 570670 257618 570906 257854
rect 570350 257298 570586 257534
rect 570670 257298 570906 257534
rect 13198 226118 13434 226354
rect 13518 226118 13754 226354
rect 13198 225798 13434 226034
rect 13518 225798 13754 226034
rect 167826 226118 168062 226354
rect 168146 226118 168382 226354
rect 167826 225798 168062 226034
rect 168146 225798 168382 226034
rect 203826 226118 204062 226354
rect 204146 226118 204382 226354
rect 203826 225798 204062 226034
rect 204146 225798 204382 226034
rect 239826 226118 240062 226354
rect 240146 226118 240382 226354
rect 239826 225798 240062 226034
rect 240146 225798 240382 226034
rect 275826 226118 276062 226354
rect 276146 226118 276382 226354
rect 275826 225798 276062 226034
rect 276146 225798 276382 226034
rect 311826 226118 312062 226354
rect 312146 226118 312382 226354
rect 311826 225798 312062 226034
rect 312146 225798 312382 226034
rect 347826 226118 348062 226354
rect 348146 226118 348382 226354
rect 347826 225798 348062 226034
rect 348146 225798 348382 226034
rect 383826 226118 384062 226354
rect 384146 226118 384382 226354
rect 383826 225798 384062 226034
rect 384146 225798 384382 226034
rect 419826 226118 420062 226354
rect 420146 226118 420382 226354
rect 419826 225798 420062 226034
rect 420146 225798 420382 226034
rect 563826 226118 564062 226354
rect 564146 226118 564382 226354
rect 563826 225798 564062 226034
rect 564146 225798 564382 226034
rect 582326 226118 582562 226354
rect 582646 226118 582882 226354
rect 582326 225798 582562 226034
rect 582646 225798 582882 226034
rect -1974 221618 -1738 221854
rect -1654 221618 -1418 221854
rect -1974 221298 -1738 221534
rect -1654 221298 -1418 221534
rect 5826 221618 6062 221854
rect 6146 221618 6382 221854
rect 5826 221298 6062 221534
rect 6146 221298 6382 221534
rect 185826 221618 186062 221854
rect 186146 221618 186382 221854
rect 185826 221298 186062 221534
rect 186146 221298 186382 221534
rect 221826 221618 222062 221854
rect 222146 221618 222382 221854
rect 221826 221298 222062 221534
rect 222146 221298 222382 221534
rect 257826 221618 258062 221854
rect 258146 221618 258382 221854
rect 257826 221298 258062 221534
rect 258146 221298 258382 221534
rect 293826 221618 294062 221854
rect 294146 221618 294382 221854
rect 293826 221298 294062 221534
rect 294146 221298 294382 221534
rect 329826 221618 330062 221854
rect 330146 221618 330382 221854
rect 329826 221298 330062 221534
rect 330146 221298 330382 221534
rect 365826 221618 366062 221854
rect 366146 221618 366382 221854
rect 365826 221298 366062 221534
rect 366146 221298 366382 221534
rect 401826 221618 402062 221854
rect 402146 221618 402382 221854
rect 401826 221298 402062 221534
rect 402146 221298 402382 221534
rect 570350 221618 570586 221854
rect 570670 221618 570906 221854
rect 570350 221298 570586 221534
rect 570670 221298 570906 221534
rect 13198 190118 13434 190354
rect 13518 190118 13754 190354
rect 13198 189798 13434 190034
rect 13518 189798 13754 190034
rect 167826 190118 168062 190354
rect 168146 190118 168382 190354
rect 167826 189798 168062 190034
rect 168146 189798 168382 190034
rect 203826 190118 204062 190354
rect 204146 190118 204382 190354
rect 203826 189798 204062 190034
rect 204146 189798 204382 190034
rect 239826 190118 240062 190354
rect 240146 190118 240382 190354
rect 239826 189798 240062 190034
rect 240146 189798 240382 190034
rect 275826 190118 276062 190354
rect 276146 190118 276382 190354
rect 275826 189798 276062 190034
rect 276146 189798 276382 190034
rect 311826 190118 312062 190354
rect 312146 190118 312382 190354
rect 311826 189798 312062 190034
rect 312146 189798 312382 190034
rect 347826 190118 348062 190354
rect 348146 190118 348382 190354
rect 347826 189798 348062 190034
rect 348146 189798 348382 190034
rect 383826 190118 384062 190354
rect 384146 190118 384382 190354
rect 383826 189798 384062 190034
rect 384146 189798 384382 190034
rect 419826 190118 420062 190354
rect 420146 190118 420382 190354
rect 419826 189798 420062 190034
rect 420146 189798 420382 190034
rect 563826 190118 564062 190354
rect 564146 190118 564382 190354
rect 563826 189798 564062 190034
rect 564146 189798 564382 190034
rect 582326 190118 582562 190354
rect 582646 190118 582882 190354
rect 582326 189798 582562 190034
rect 582646 189798 582882 190034
rect -1974 185618 -1738 185854
rect -1654 185618 -1418 185854
rect -1974 185298 -1738 185534
rect -1654 185298 -1418 185534
rect 5826 185618 6062 185854
rect 6146 185618 6382 185854
rect 5826 185298 6062 185534
rect 6146 185298 6382 185534
rect 185826 185618 186062 185854
rect 186146 185618 186382 185854
rect 185826 185298 186062 185534
rect 186146 185298 186382 185534
rect 221826 185618 222062 185854
rect 222146 185618 222382 185854
rect 221826 185298 222062 185534
rect 222146 185298 222382 185534
rect 257826 185618 258062 185854
rect 258146 185618 258382 185854
rect 257826 185298 258062 185534
rect 258146 185298 258382 185534
rect 293826 185618 294062 185854
rect 294146 185618 294382 185854
rect 293826 185298 294062 185534
rect 294146 185298 294382 185534
rect 329826 185618 330062 185854
rect 330146 185618 330382 185854
rect 329826 185298 330062 185534
rect 330146 185298 330382 185534
rect 365826 185618 366062 185854
rect 366146 185618 366382 185854
rect 365826 185298 366062 185534
rect 366146 185298 366382 185534
rect 401826 185618 402062 185854
rect 402146 185618 402382 185854
rect 401826 185298 402062 185534
rect 402146 185298 402382 185534
rect 570350 185618 570586 185854
rect 570670 185618 570906 185854
rect 570350 185298 570586 185534
rect 570670 185298 570906 185534
rect 13198 154118 13434 154354
rect 13518 154118 13754 154354
rect 13198 153798 13434 154034
rect 13518 153798 13754 154034
rect 167826 154118 168062 154354
rect 168146 154118 168382 154354
rect 167826 153798 168062 154034
rect 168146 153798 168382 154034
rect 203826 154118 204062 154354
rect 204146 154118 204382 154354
rect 203826 153798 204062 154034
rect 204146 153798 204382 154034
rect 239826 154118 240062 154354
rect 240146 154118 240382 154354
rect 239826 153798 240062 154034
rect 240146 153798 240382 154034
rect 275826 154118 276062 154354
rect 276146 154118 276382 154354
rect 275826 153798 276062 154034
rect 276146 153798 276382 154034
rect 311826 154118 312062 154354
rect 312146 154118 312382 154354
rect 311826 153798 312062 154034
rect 312146 153798 312382 154034
rect 347826 154118 348062 154354
rect 348146 154118 348382 154354
rect 347826 153798 348062 154034
rect 348146 153798 348382 154034
rect 383826 154118 384062 154354
rect 384146 154118 384382 154354
rect 383826 153798 384062 154034
rect 384146 153798 384382 154034
rect 419826 154118 420062 154354
rect 420146 154118 420382 154354
rect 419826 153798 420062 154034
rect 420146 153798 420382 154034
rect 563826 154118 564062 154354
rect 564146 154118 564382 154354
rect 563826 153798 564062 154034
rect 564146 153798 564382 154034
rect 582326 154118 582562 154354
rect 582646 154118 582882 154354
rect 582326 153798 582562 154034
rect 582646 153798 582882 154034
rect -1974 149618 -1738 149854
rect -1654 149618 -1418 149854
rect -1974 149298 -1738 149534
rect -1654 149298 -1418 149534
rect 5826 149618 6062 149854
rect 6146 149618 6382 149854
rect 5826 149298 6062 149534
rect 6146 149298 6382 149534
rect 185826 149618 186062 149854
rect 186146 149618 186382 149854
rect 185826 149298 186062 149534
rect 186146 149298 186382 149534
rect 221826 149618 222062 149854
rect 222146 149618 222382 149854
rect 221826 149298 222062 149534
rect 222146 149298 222382 149534
rect 257826 149618 258062 149854
rect 258146 149618 258382 149854
rect 257826 149298 258062 149534
rect 258146 149298 258382 149534
rect 293826 149618 294062 149854
rect 294146 149618 294382 149854
rect 293826 149298 294062 149534
rect 294146 149298 294382 149534
rect 329826 149618 330062 149854
rect 330146 149618 330382 149854
rect 329826 149298 330062 149534
rect 330146 149298 330382 149534
rect 365826 149618 366062 149854
rect 366146 149618 366382 149854
rect 365826 149298 366062 149534
rect 366146 149298 366382 149534
rect 401826 149618 402062 149854
rect 402146 149618 402382 149854
rect 401826 149298 402062 149534
rect 402146 149298 402382 149534
rect 570350 149618 570586 149854
rect 570670 149618 570906 149854
rect 570350 149298 570586 149534
rect 570670 149298 570906 149534
rect 13198 118118 13434 118354
rect 13518 118118 13754 118354
rect 13198 117798 13434 118034
rect 13518 117798 13754 118034
rect 167826 118118 168062 118354
rect 168146 118118 168382 118354
rect 167826 117798 168062 118034
rect 168146 117798 168382 118034
rect 203826 118118 204062 118354
rect 204146 118118 204382 118354
rect 203826 117798 204062 118034
rect 204146 117798 204382 118034
rect 239826 118118 240062 118354
rect 240146 118118 240382 118354
rect 239826 117798 240062 118034
rect 240146 117798 240382 118034
rect 275826 118118 276062 118354
rect 276146 118118 276382 118354
rect 275826 117798 276062 118034
rect 276146 117798 276382 118034
rect 311826 118118 312062 118354
rect 312146 118118 312382 118354
rect 311826 117798 312062 118034
rect 312146 117798 312382 118034
rect 347826 118118 348062 118354
rect 348146 118118 348382 118354
rect 347826 117798 348062 118034
rect 348146 117798 348382 118034
rect 383826 118118 384062 118354
rect 384146 118118 384382 118354
rect 383826 117798 384062 118034
rect 384146 117798 384382 118034
rect 419826 118118 420062 118354
rect 420146 118118 420382 118354
rect 419826 117798 420062 118034
rect 420146 117798 420382 118034
rect 563826 118118 564062 118354
rect 564146 118118 564382 118354
rect 563826 117798 564062 118034
rect 564146 117798 564382 118034
rect 582326 118118 582562 118354
rect 582646 118118 582882 118354
rect 582326 117798 582562 118034
rect 582646 117798 582882 118034
rect -1974 113618 -1738 113854
rect -1654 113618 -1418 113854
rect -1974 113298 -1738 113534
rect -1654 113298 -1418 113534
rect 5826 113618 6062 113854
rect 6146 113618 6382 113854
rect 5826 113298 6062 113534
rect 6146 113298 6382 113534
rect 173094 113618 173330 113854
rect 173414 113618 173650 113854
rect 173094 113298 173330 113534
rect 173414 113298 173650 113534
rect 293826 113618 294062 113854
rect 294146 113618 294382 113854
rect 293826 113298 294062 113534
rect 294146 113298 294382 113534
rect 401826 113618 402062 113854
rect 402146 113618 402382 113854
rect 401826 113298 402062 113534
rect 402146 113298 402382 113534
rect 570350 113618 570586 113854
rect 570670 113618 570906 113854
rect 570350 113298 570586 113534
rect 570670 113298 570906 113534
rect 13198 82118 13434 82354
rect 13518 82118 13754 82354
rect 13198 81798 13434 82034
rect 13518 81798 13754 82034
rect 167826 82118 168062 82354
rect 168146 82118 168382 82354
rect 167826 81798 168062 82034
rect 168146 81798 168382 82034
rect 291590 82118 291826 82354
rect 291910 82118 292146 82354
rect 291590 81798 291826 82034
rect 291910 81798 292146 82034
rect 419826 82118 420062 82354
rect 420146 82118 420382 82354
rect 419826 81798 420062 82034
rect 420146 81798 420382 82034
rect 563826 82118 564062 82354
rect 564146 82118 564382 82354
rect 563826 81798 564062 82034
rect 564146 81798 564382 82034
rect 582326 82118 582562 82354
rect 582646 82118 582882 82354
rect 582326 81798 582562 82034
rect 582646 81798 582882 82034
rect -1974 77618 -1738 77854
rect -1654 77618 -1418 77854
rect -1974 77298 -1738 77534
rect -1654 77298 -1418 77534
rect 5826 77618 6062 77854
rect 6146 77618 6382 77854
rect 5826 77298 6062 77534
rect 6146 77298 6382 77534
rect 173094 77618 173330 77854
rect 173414 77618 173650 77854
rect 173094 77298 173330 77534
rect 173414 77298 173650 77534
rect 293826 77618 294062 77854
rect 294146 77618 294382 77854
rect 293826 77298 294062 77534
rect 294146 77298 294382 77534
rect 401826 77618 402062 77854
rect 402146 77618 402382 77854
rect 401826 77298 402062 77534
rect 402146 77298 402382 77534
rect 570350 77618 570586 77854
rect 570670 77618 570906 77854
rect 570350 77298 570586 77534
rect 570670 77298 570906 77534
rect 13198 46118 13434 46354
rect 13518 46118 13754 46354
rect 13198 45798 13434 46034
rect 13518 45798 13754 46034
rect 167826 46118 168062 46354
rect 168146 46118 168382 46354
rect 167826 45798 168062 46034
rect 168146 45798 168382 46034
rect 291590 46118 291826 46354
rect 291910 46118 292146 46354
rect 291590 45798 291826 46034
rect 291910 45798 292146 46034
rect 419826 46118 420062 46354
rect 420146 46118 420382 46354
rect 419826 45798 420062 46034
rect 420146 45798 420382 46034
rect 563826 46118 564062 46354
rect 564146 46118 564382 46354
rect 563826 45798 564062 46034
rect 564146 45798 564382 46034
rect 582326 46118 582562 46354
rect 582646 46118 582882 46354
rect 582326 45798 582562 46034
rect 582646 45798 582882 46034
rect -1974 41618 -1738 41854
rect -1654 41618 -1418 41854
rect -1974 41298 -1738 41534
rect -1654 41298 -1418 41534
rect 5826 41618 6062 41854
rect 6146 41618 6382 41854
rect 5826 41298 6062 41534
rect 6146 41298 6382 41534
rect 173094 41618 173330 41854
rect 173414 41618 173650 41854
rect 173094 41298 173330 41534
rect 173414 41298 173650 41534
rect 293826 41618 294062 41854
rect 294146 41618 294382 41854
rect 293826 41298 294062 41534
rect 294146 41298 294382 41534
rect 401826 41618 402062 41854
rect 402146 41618 402382 41854
rect 401826 41298 402062 41534
rect 402146 41298 402382 41534
rect 570350 41618 570586 41854
rect 570670 41618 570906 41854
rect 570350 41298 570586 41534
rect 570670 41298 570906 41534
rect 23826 10118 24062 10354
rect 24146 10118 24382 10354
rect 23826 9798 24062 10034
rect 24146 9798 24382 10034
rect 59826 10118 60062 10354
rect 60146 10118 60382 10354
rect 59826 9798 60062 10034
rect 60146 9798 60382 10034
rect 95826 10118 96062 10354
rect 96146 10118 96382 10354
rect 95826 9798 96062 10034
rect 96146 9798 96382 10034
rect 131826 10118 132062 10354
rect 132146 10118 132382 10354
rect 131826 9798 132062 10034
rect 132146 9798 132382 10034
rect 167826 10118 168062 10354
rect 168146 10118 168382 10354
rect 167826 9798 168062 10034
rect 168146 9798 168382 10034
rect 203826 10118 204062 10354
rect 204146 10118 204382 10354
rect 203826 9798 204062 10034
rect 204146 9798 204382 10034
rect 239826 10118 240062 10354
rect 240146 10118 240382 10354
rect 239826 9798 240062 10034
rect 240146 9798 240382 10034
rect 275826 10118 276062 10354
rect 276146 10118 276382 10354
rect 275826 9798 276062 10034
rect 276146 9798 276382 10034
rect 311826 10118 312062 10354
rect 312146 10118 312382 10354
rect 311826 9798 312062 10034
rect 312146 9798 312382 10034
rect 347826 10118 348062 10354
rect 348146 10118 348382 10354
rect 347826 9798 348062 10034
rect 348146 9798 348382 10034
rect 383826 10118 384062 10354
rect 384146 10118 384382 10354
rect 383826 9798 384062 10034
rect 384146 9798 384382 10034
rect 419826 10118 420062 10354
rect 420146 10118 420382 10354
rect 419826 9798 420062 10034
rect 420146 9798 420382 10034
rect 455826 10118 456062 10354
rect 456146 10118 456382 10354
rect 455826 9798 456062 10034
rect 456146 9798 456382 10034
rect 491826 10118 492062 10354
rect 492146 10118 492382 10354
rect 491826 9798 492062 10034
rect 492146 9798 492382 10034
rect 527826 10118 528062 10354
rect 528146 10118 528382 10354
rect 527826 9798 528062 10034
rect 528146 9798 528382 10034
rect 563826 10118 564062 10354
rect 564146 10118 564382 10354
rect 563826 9798 564062 10034
rect 564146 9798 564382 10034
rect 582326 10118 582562 10354
rect 582646 10118 582882 10354
rect 582326 9798 582562 10034
rect 582646 9798 582882 10034
rect -1974 5618 -1738 5854
rect -1654 5618 -1418 5854
rect -1974 5298 -1738 5534
rect -1654 5298 -1418 5534
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 689618 585578 689854
rect 585662 689618 585898 689854
rect 585342 689298 585578 689534
rect 585662 689298 585898 689534
rect 585342 653618 585578 653854
rect 585662 653618 585898 653854
rect 585342 653298 585578 653534
rect 585662 653298 585898 653534
rect 585342 617618 585578 617854
rect 585662 617618 585898 617854
rect 585342 617298 585578 617534
rect 585662 617298 585898 617534
rect 585342 581618 585578 581854
rect 585662 581618 585898 581854
rect 585342 581298 585578 581534
rect 585662 581298 585898 581534
rect 585342 545618 585578 545854
rect 585662 545618 585898 545854
rect 585342 545298 585578 545534
rect 585662 545298 585898 545534
rect 585342 509618 585578 509854
rect 585662 509618 585898 509854
rect 585342 509298 585578 509534
rect 585662 509298 585898 509534
rect 585342 473618 585578 473854
rect 585662 473618 585898 473854
rect 585342 473298 585578 473534
rect 585662 473298 585898 473534
rect 585342 437618 585578 437854
rect 585662 437618 585898 437854
rect 585342 437298 585578 437534
rect 585662 437298 585898 437534
rect 585342 401618 585578 401854
rect 585662 401618 585898 401854
rect 585342 401298 585578 401534
rect 585662 401298 585898 401534
rect 585342 365618 585578 365854
rect 585662 365618 585898 365854
rect 585342 365298 585578 365534
rect 585662 365298 585898 365534
rect 585342 329618 585578 329854
rect 585662 329618 585898 329854
rect 585342 329298 585578 329534
rect 585662 329298 585898 329534
rect 585342 293618 585578 293854
rect 585662 293618 585898 293854
rect 585342 293298 585578 293534
rect 585662 293298 585898 293534
rect 585342 257618 585578 257854
rect 585662 257618 585898 257854
rect 585342 257298 585578 257534
rect 585662 257298 585898 257534
rect 585342 221618 585578 221854
rect 585662 221618 585898 221854
rect 585342 221298 585578 221534
rect 585662 221298 585898 221534
rect 585342 185618 585578 185854
rect 585662 185618 585898 185854
rect 585342 185298 585578 185534
rect 585662 185298 585898 185534
rect 585342 149618 585578 149854
rect 585662 149618 585898 149854
rect 585342 149298 585578 149534
rect 585662 149298 585898 149534
rect 585342 113618 585578 113854
rect 585662 113618 585898 113854
rect 585342 113298 585578 113534
rect 585662 113298 585898 113534
rect 585342 77618 585578 77854
rect 585662 77618 585898 77854
rect 585342 77298 585578 77534
rect 585662 77298 585898 77534
rect 585342 41618 585578 41854
rect 585662 41618 585898 41854
rect 585342 41298 585578 41534
rect 585662 41298 585898 41534
rect 585342 5618 585578 5854
rect 585662 5618 585898 5854
rect 585342 5298 585578 5534
rect 585662 5298 585898 5534
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 694118 586538 694354
rect 586622 694118 586858 694354
rect 586302 693798 586538 694034
rect 586622 693798 586858 694034
rect 586302 658118 586538 658354
rect 586622 658118 586858 658354
rect 586302 657798 586538 658034
rect 586622 657798 586858 658034
rect 586302 622118 586538 622354
rect 586622 622118 586858 622354
rect 586302 621798 586538 622034
rect 586622 621798 586858 622034
rect 586302 586118 586538 586354
rect 586622 586118 586858 586354
rect 586302 585798 586538 586034
rect 586622 585798 586858 586034
rect 586302 550118 586538 550354
rect 586622 550118 586858 550354
rect 586302 549798 586538 550034
rect 586622 549798 586858 550034
rect 586302 514118 586538 514354
rect 586622 514118 586858 514354
rect 586302 513798 586538 514034
rect 586622 513798 586858 514034
rect 586302 478118 586538 478354
rect 586622 478118 586858 478354
rect 586302 477798 586538 478034
rect 586622 477798 586858 478034
rect 586302 442118 586538 442354
rect 586622 442118 586858 442354
rect 586302 441798 586538 442034
rect 586622 441798 586858 442034
rect 586302 406118 586538 406354
rect 586622 406118 586858 406354
rect 586302 405798 586538 406034
rect 586622 405798 586858 406034
rect 586302 370118 586538 370354
rect 586622 370118 586858 370354
rect 586302 369798 586538 370034
rect 586622 369798 586858 370034
rect 586302 334118 586538 334354
rect 586622 334118 586858 334354
rect 586302 333798 586538 334034
rect 586622 333798 586858 334034
rect 586302 298118 586538 298354
rect 586622 298118 586858 298354
rect 586302 297798 586538 298034
rect 586622 297798 586858 298034
rect 586302 262118 586538 262354
rect 586622 262118 586858 262354
rect 586302 261798 586538 262034
rect 586622 261798 586858 262034
rect 586302 226118 586538 226354
rect 586622 226118 586858 226354
rect 586302 225798 586538 226034
rect 586622 225798 586858 226034
rect 586302 190118 586538 190354
rect 586622 190118 586858 190354
rect 586302 189798 586538 190034
rect 586622 189798 586858 190034
rect 586302 154118 586538 154354
rect 586622 154118 586858 154354
rect 586302 153798 586538 154034
rect 586622 153798 586858 154034
rect 586302 118118 586538 118354
rect 586622 118118 586858 118354
rect 586302 117798 586538 118034
rect 586622 117798 586858 118034
rect 586302 82118 586538 82354
rect 586622 82118 586858 82354
rect 586302 81798 586538 82034
rect 586622 81798 586858 82034
rect 586302 46118 586538 46354
rect 586622 46118 586858 46354
rect 586302 45798 586538 46034
rect 586622 45798 586858 46034
rect 586302 10118 586538 10354
rect 586622 10118 586858 10354
rect 586302 9798 586538 10034
rect 586622 9798 586858 10034
rect 582326 -1542 582562 -1306
rect 582646 -1542 582882 -1306
rect 582326 -1862 582562 -1626
rect 582646 -1862 582882 -1626
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 582326 705798
rect 582562 705562 582646 705798
rect 582882 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 582326 705478
rect 582562 705242 582646 705478
rect 582882 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 694354 592650 694386
rect -8726 694118 -2934 694354
rect -2698 694118 -2614 694354
rect -2378 694118 23826 694354
rect 24062 694118 24146 694354
rect 24382 694118 59826 694354
rect 60062 694118 60146 694354
rect 60382 694118 95826 694354
rect 96062 694118 96146 694354
rect 96382 694118 131826 694354
rect 132062 694118 132146 694354
rect 132382 694118 167826 694354
rect 168062 694118 168146 694354
rect 168382 694118 203826 694354
rect 204062 694118 204146 694354
rect 204382 694118 239826 694354
rect 240062 694118 240146 694354
rect 240382 694118 275826 694354
rect 276062 694118 276146 694354
rect 276382 694118 311826 694354
rect 312062 694118 312146 694354
rect 312382 694118 347826 694354
rect 348062 694118 348146 694354
rect 348382 694118 383826 694354
rect 384062 694118 384146 694354
rect 384382 694118 419826 694354
rect 420062 694118 420146 694354
rect 420382 694118 455826 694354
rect 456062 694118 456146 694354
rect 456382 694118 491826 694354
rect 492062 694118 492146 694354
rect 492382 694118 527826 694354
rect 528062 694118 528146 694354
rect 528382 694118 563826 694354
rect 564062 694118 564146 694354
rect 564382 694118 582326 694354
rect 582562 694118 582646 694354
rect 582882 694118 586302 694354
rect 586538 694118 586622 694354
rect 586858 694118 592650 694354
rect -8726 694034 592650 694118
rect -8726 693798 -2934 694034
rect -2698 693798 -2614 694034
rect -2378 693798 23826 694034
rect 24062 693798 24146 694034
rect 24382 693798 59826 694034
rect 60062 693798 60146 694034
rect 60382 693798 95826 694034
rect 96062 693798 96146 694034
rect 96382 693798 131826 694034
rect 132062 693798 132146 694034
rect 132382 693798 167826 694034
rect 168062 693798 168146 694034
rect 168382 693798 203826 694034
rect 204062 693798 204146 694034
rect 204382 693798 239826 694034
rect 240062 693798 240146 694034
rect 240382 693798 275826 694034
rect 276062 693798 276146 694034
rect 276382 693798 311826 694034
rect 312062 693798 312146 694034
rect 312382 693798 347826 694034
rect 348062 693798 348146 694034
rect 348382 693798 383826 694034
rect 384062 693798 384146 694034
rect 384382 693798 419826 694034
rect 420062 693798 420146 694034
rect 420382 693798 455826 694034
rect 456062 693798 456146 694034
rect 456382 693798 491826 694034
rect 492062 693798 492146 694034
rect 492382 693798 527826 694034
rect 528062 693798 528146 694034
rect 528382 693798 563826 694034
rect 564062 693798 564146 694034
rect 564382 693798 582326 694034
rect 582562 693798 582646 694034
rect 582882 693798 586302 694034
rect 586538 693798 586622 694034
rect 586858 693798 592650 694034
rect -8726 693766 592650 693798
rect -8726 689854 592650 689886
rect -8726 689618 -1974 689854
rect -1738 689618 -1654 689854
rect -1418 689618 5826 689854
rect 6062 689618 6146 689854
rect 6382 689618 41826 689854
rect 42062 689618 42146 689854
rect 42382 689618 77826 689854
rect 78062 689618 78146 689854
rect 78382 689618 113826 689854
rect 114062 689618 114146 689854
rect 114382 689618 149826 689854
rect 150062 689618 150146 689854
rect 150382 689618 185826 689854
rect 186062 689618 186146 689854
rect 186382 689618 221826 689854
rect 222062 689618 222146 689854
rect 222382 689618 257826 689854
rect 258062 689618 258146 689854
rect 258382 689618 293826 689854
rect 294062 689618 294146 689854
rect 294382 689618 329826 689854
rect 330062 689618 330146 689854
rect 330382 689618 365826 689854
rect 366062 689618 366146 689854
rect 366382 689618 401826 689854
rect 402062 689618 402146 689854
rect 402382 689618 437826 689854
rect 438062 689618 438146 689854
rect 438382 689618 473826 689854
rect 474062 689618 474146 689854
rect 474382 689618 509826 689854
rect 510062 689618 510146 689854
rect 510382 689618 545826 689854
rect 546062 689618 546146 689854
rect 546382 689618 585342 689854
rect 585578 689618 585662 689854
rect 585898 689618 592650 689854
rect -8726 689534 592650 689618
rect -8726 689298 -1974 689534
rect -1738 689298 -1654 689534
rect -1418 689298 5826 689534
rect 6062 689298 6146 689534
rect 6382 689298 41826 689534
rect 42062 689298 42146 689534
rect 42382 689298 77826 689534
rect 78062 689298 78146 689534
rect 78382 689298 113826 689534
rect 114062 689298 114146 689534
rect 114382 689298 149826 689534
rect 150062 689298 150146 689534
rect 150382 689298 185826 689534
rect 186062 689298 186146 689534
rect 186382 689298 221826 689534
rect 222062 689298 222146 689534
rect 222382 689298 257826 689534
rect 258062 689298 258146 689534
rect 258382 689298 293826 689534
rect 294062 689298 294146 689534
rect 294382 689298 329826 689534
rect 330062 689298 330146 689534
rect 330382 689298 365826 689534
rect 366062 689298 366146 689534
rect 366382 689298 401826 689534
rect 402062 689298 402146 689534
rect 402382 689298 437826 689534
rect 438062 689298 438146 689534
rect 438382 689298 473826 689534
rect 474062 689298 474146 689534
rect 474382 689298 509826 689534
rect 510062 689298 510146 689534
rect 510382 689298 545826 689534
rect 546062 689298 546146 689534
rect 546382 689298 585342 689534
rect 585578 689298 585662 689534
rect 585898 689298 592650 689534
rect -8726 689266 592650 689298
rect -8726 658354 592650 658386
rect -8726 658118 -2934 658354
rect -2698 658118 -2614 658354
rect -2378 658118 13198 658354
rect 13434 658118 13518 658354
rect 13754 658118 167826 658354
rect 168062 658118 168146 658354
rect 168382 658118 291590 658354
rect 291826 658118 291910 658354
rect 292146 658118 419826 658354
rect 420062 658118 420146 658354
rect 420382 658118 563826 658354
rect 564062 658118 564146 658354
rect 564382 658118 582326 658354
rect 582562 658118 582646 658354
rect 582882 658118 586302 658354
rect 586538 658118 586622 658354
rect 586858 658118 592650 658354
rect -8726 658034 592650 658118
rect -8726 657798 -2934 658034
rect -2698 657798 -2614 658034
rect -2378 657798 13198 658034
rect 13434 657798 13518 658034
rect 13754 657798 167826 658034
rect 168062 657798 168146 658034
rect 168382 657798 291590 658034
rect 291826 657798 291910 658034
rect 292146 657798 419826 658034
rect 420062 657798 420146 658034
rect 420382 657798 563826 658034
rect 564062 657798 564146 658034
rect 564382 657798 582326 658034
rect 582562 657798 582646 658034
rect 582882 657798 586302 658034
rect 586538 657798 586622 658034
rect 586858 657798 592650 658034
rect -8726 657766 592650 657798
rect -8726 653854 592650 653886
rect -8726 653618 -1974 653854
rect -1738 653618 -1654 653854
rect -1418 653618 5826 653854
rect 6062 653618 6146 653854
rect 6382 653618 173094 653854
rect 173330 653618 173414 653854
rect 173650 653618 293826 653854
rect 294062 653618 294146 653854
rect 294382 653618 401826 653854
rect 402062 653618 402146 653854
rect 402382 653618 570350 653854
rect 570586 653618 570670 653854
rect 570906 653618 585342 653854
rect 585578 653618 585662 653854
rect 585898 653618 592650 653854
rect -8726 653534 592650 653618
rect -8726 653298 -1974 653534
rect -1738 653298 -1654 653534
rect -1418 653298 5826 653534
rect 6062 653298 6146 653534
rect 6382 653298 173094 653534
rect 173330 653298 173414 653534
rect 173650 653298 293826 653534
rect 294062 653298 294146 653534
rect 294382 653298 401826 653534
rect 402062 653298 402146 653534
rect 402382 653298 570350 653534
rect 570586 653298 570670 653534
rect 570906 653298 585342 653534
rect 585578 653298 585662 653534
rect 585898 653298 592650 653534
rect -8726 653266 592650 653298
rect -8726 622354 592650 622386
rect -8726 622118 -2934 622354
rect -2698 622118 -2614 622354
rect -2378 622118 13198 622354
rect 13434 622118 13518 622354
rect 13754 622118 167826 622354
rect 168062 622118 168146 622354
rect 168382 622118 291590 622354
rect 291826 622118 291910 622354
rect 292146 622118 419826 622354
rect 420062 622118 420146 622354
rect 420382 622118 563826 622354
rect 564062 622118 564146 622354
rect 564382 622118 582326 622354
rect 582562 622118 582646 622354
rect 582882 622118 586302 622354
rect 586538 622118 586622 622354
rect 586858 622118 592650 622354
rect -8726 622034 592650 622118
rect -8726 621798 -2934 622034
rect -2698 621798 -2614 622034
rect -2378 621798 13198 622034
rect 13434 621798 13518 622034
rect 13754 621798 167826 622034
rect 168062 621798 168146 622034
rect 168382 621798 291590 622034
rect 291826 621798 291910 622034
rect 292146 621798 419826 622034
rect 420062 621798 420146 622034
rect 420382 621798 563826 622034
rect 564062 621798 564146 622034
rect 564382 621798 582326 622034
rect 582562 621798 582646 622034
rect 582882 621798 586302 622034
rect 586538 621798 586622 622034
rect 586858 621798 592650 622034
rect -8726 621766 592650 621798
rect -8726 617854 592650 617886
rect -8726 617618 -1974 617854
rect -1738 617618 -1654 617854
rect -1418 617618 5826 617854
rect 6062 617618 6146 617854
rect 6382 617618 173094 617854
rect 173330 617618 173414 617854
rect 173650 617618 293826 617854
rect 294062 617618 294146 617854
rect 294382 617618 401826 617854
rect 402062 617618 402146 617854
rect 402382 617618 570350 617854
rect 570586 617618 570670 617854
rect 570906 617618 585342 617854
rect 585578 617618 585662 617854
rect 585898 617618 592650 617854
rect -8726 617534 592650 617618
rect -8726 617298 -1974 617534
rect -1738 617298 -1654 617534
rect -1418 617298 5826 617534
rect 6062 617298 6146 617534
rect 6382 617298 173094 617534
rect 173330 617298 173414 617534
rect 173650 617298 293826 617534
rect 294062 617298 294146 617534
rect 294382 617298 401826 617534
rect 402062 617298 402146 617534
rect 402382 617298 570350 617534
rect 570586 617298 570670 617534
rect 570906 617298 585342 617534
rect 585578 617298 585662 617534
rect 585898 617298 592650 617534
rect -8726 617266 592650 617298
rect -8726 586354 592650 586386
rect -8726 586118 -2934 586354
rect -2698 586118 -2614 586354
rect -2378 586118 23826 586354
rect 24062 586118 24146 586354
rect 24382 586118 59826 586354
rect 60062 586118 60146 586354
rect 60382 586118 95826 586354
rect 96062 586118 96146 586354
rect 96382 586118 131826 586354
rect 132062 586118 132146 586354
rect 132382 586118 167826 586354
rect 168062 586118 168146 586354
rect 168382 586118 203826 586354
rect 204062 586118 204146 586354
rect 204382 586118 239826 586354
rect 240062 586118 240146 586354
rect 240382 586118 275826 586354
rect 276062 586118 276146 586354
rect 276382 586118 311826 586354
rect 312062 586118 312146 586354
rect 312382 586118 347826 586354
rect 348062 586118 348146 586354
rect 348382 586118 383826 586354
rect 384062 586118 384146 586354
rect 384382 586118 419826 586354
rect 420062 586118 420146 586354
rect 420382 586118 455826 586354
rect 456062 586118 456146 586354
rect 456382 586118 491826 586354
rect 492062 586118 492146 586354
rect 492382 586118 527826 586354
rect 528062 586118 528146 586354
rect 528382 586118 563826 586354
rect 564062 586118 564146 586354
rect 564382 586118 582326 586354
rect 582562 586118 582646 586354
rect 582882 586118 586302 586354
rect 586538 586118 586622 586354
rect 586858 586118 592650 586354
rect -8726 586034 592650 586118
rect -8726 585798 -2934 586034
rect -2698 585798 -2614 586034
rect -2378 585798 23826 586034
rect 24062 585798 24146 586034
rect 24382 585798 59826 586034
rect 60062 585798 60146 586034
rect 60382 585798 95826 586034
rect 96062 585798 96146 586034
rect 96382 585798 131826 586034
rect 132062 585798 132146 586034
rect 132382 585798 167826 586034
rect 168062 585798 168146 586034
rect 168382 585798 203826 586034
rect 204062 585798 204146 586034
rect 204382 585798 239826 586034
rect 240062 585798 240146 586034
rect 240382 585798 275826 586034
rect 276062 585798 276146 586034
rect 276382 585798 311826 586034
rect 312062 585798 312146 586034
rect 312382 585798 347826 586034
rect 348062 585798 348146 586034
rect 348382 585798 383826 586034
rect 384062 585798 384146 586034
rect 384382 585798 419826 586034
rect 420062 585798 420146 586034
rect 420382 585798 455826 586034
rect 456062 585798 456146 586034
rect 456382 585798 491826 586034
rect 492062 585798 492146 586034
rect 492382 585798 527826 586034
rect 528062 585798 528146 586034
rect 528382 585798 563826 586034
rect 564062 585798 564146 586034
rect 564382 585798 582326 586034
rect 582562 585798 582646 586034
rect 582882 585798 586302 586034
rect 586538 585798 586622 586034
rect 586858 585798 592650 586034
rect -8726 585766 592650 585798
rect -8726 581854 592650 581886
rect -8726 581618 -1974 581854
rect -1738 581618 -1654 581854
rect -1418 581618 5826 581854
rect 6062 581618 6146 581854
rect 6382 581618 41826 581854
rect 42062 581618 42146 581854
rect 42382 581618 77826 581854
rect 78062 581618 78146 581854
rect 78382 581618 113826 581854
rect 114062 581618 114146 581854
rect 114382 581618 149826 581854
rect 150062 581618 150146 581854
rect 150382 581618 185826 581854
rect 186062 581618 186146 581854
rect 186382 581618 221826 581854
rect 222062 581618 222146 581854
rect 222382 581618 257826 581854
rect 258062 581618 258146 581854
rect 258382 581618 293826 581854
rect 294062 581618 294146 581854
rect 294382 581618 329826 581854
rect 330062 581618 330146 581854
rect 330382 581618 365826 581854
rect 366062 581618 366146 581854
rect 366382 581618 401826 581854
rect 402062 581618 402146 581854
rect 402382 581618 437826 581854
rect 438062 581618 438146 581854
rect 438382 581618 473826 581854
rect 474062 581618 474146 581854
rect 474382 581618 509826 581854
rect 510062 581618 510146 581854
rect 510382 581618 545826 581854
rect 546062 581618 546146 581854
rect 546382 581618 585342 581854
rect 585578 581618 585662 581854
rect 585898 581618 592650 581854
rect -8726 581534 592650 581618
rect -8726 581298 -1974 581534
rect -1738 581298 -1654 581534
rect -1418 581298 5826 581534
rect 6062 581298 6146 581534
rect 6382 581298 41826 581534
rect 42062 581298 42146 581534
rect 42382 581298 77826 581534
rect 78062 581298 78146 581534
rect 78382 581298 113826 581534
rect 114062 581298 114146 581534
rect 114382 581298 149826 581534
rect 150062 581298 150146 581534
rect 150382 581298 185826 581534
rect 186062 581298 186146 581534
rect 186382 581298 221826 581534
rect 222062 581298 222146 581534
rect 222382 581298 257826 581534
rect 258062 581298 258146 581534
rect 258382 581298 293826 581534
rect 294062 581298 294146 581534
rect 294382 581298 329826 581534
rect 330062 581298 330146 581534
rect 330382 581298 365826 581534
rect 366062 581298 366146 581534
rect 366382 581298 401826 581534
rect 402062 581298 402146 581534
rect 402382 581298 437826 581534
rect 438062 581298 438146 581534
rect 438382 581298 473826 581534
rect 474062 581298 474146 581534
rect 474382 581298 509826 581534
rect 510062 581298 510146 581534
rect 510382 581298 545826 581534
rect 546062 581298 546146 581534
rect 546382 581298 585342 581534
rect 585578 581298 585662 581534
rect 585898 581298 592650 581534
rect -8726 581266 592650 581298
rect -8726 550354 592650 550386
rect -8726 550118 -2934 550354
rect -2698 550118 -2614 550354
rect -2378 550118 13198 550354
rect 13434 550118 13518 550354
rect 13754 550118 167826 550354
rect 168062 550118 168146 550354
rect 168382 550118 203826 550354
rect 204062 550118 204146 550354
rect 204382 550118 239826 550354
rect 240062 550118 240146 550354
rect 240382 550118 275826 550354
rect 276062 550118 276146 550354
rect 276382 550118 311826 550354
rect 312062 550118 312146 550354
rect 312382 550118 347826 550354
rect 348062 550118 348146 550354
rect 348382 550118 383826 550354
rect 384062 550118 384146 550354
rect 384382 550118 419826 550354
rect 420062 550118 420146 550354
rect 420382 550118 563826 550354
rect 564062 550118 564146 550354
rect 564382 550118 582326 550354
rect 582562 550118 582646 550354
rect 582882 550118 586302 550354
rect 586538 550118 586622 550354
rect 586858 550118 592650 550354
rect -8726 550034 592650 550118
rect -8726 549798 -2934 550034
rect -2698 549798 -2614 550034
rect -2378 549798 13198 550034
rect 13434 549798 13518 550034
rect 13754 549798 167826 550034
rect 168062 549798 168146 550034
rect 168382 549798 203826 550034
rect 204062 549798 204146 550034
rect 204382 549798 239826 550034
rect 240062 549798 240146 550034
rect 240382 549798 275826 550034
rect 276062 549798 276146 550034
rect 276382 549798 311826 550034
rect 312062 549798 312146 550034
rect 312382 549798 347826 550034
rect 348062 549798 348146 550034
rect 348382 549798 383826 550034
rect 384062 549798 384146 550034
rect 384382 549798 419826 550034
rect 420062 549798 420146 550034
rect 420382 549798 563826 550034
rect 564062 549798 564146 550034
rect 564382 549798 582326 550034
rect 582562 549798 582646 550034
rect 582882 549798 586302 550034
rect 586538 549798 586622 550034
rect 586858 549798 592650 550034
rect -8726 549766 592650 549798
rect -8726 545854 592650 545886
rect -8726 545618 -1974 545854
rect -1738 545618 -1654 545854
rect -1418 545618 5826 545854
rect 6062 545618 6146 545854
rect 6382 545618 185826 545854
rect 186062 545618 186146 545854
rect 186382 545618 221826 545854
rect 222062 545618 222146 545854
rect 222382 545618 257826 545854
rect 258062 545618 258146 545854
rect 258382 545618 293826 545854
rect 294062 545618 294146 545854
rect 294382 545618 329826 545854
rect 330062 545618 330146 545854
rect 330382 545618 365826 545854
rect 366062 545618 366146 545854
rect 366382 545618 401826 545854
rect 402062 545618 402146 545854
rect 402382 545618 570350 545854
rect 570586 545618 570670 545854
rect 570906 545618 585342 545854
rect 585578 545618 585662 545854
rect 585898 545618 592650 545854
rect -8726 545534 592650 545618
rect -8726 545298 -1974 545534
rect -1738 545298 -1654 545534
rect -1418 545298 5826 545534
rect 6062 545298 6146 545534
rect 6382 545298 185826 545534
rect 186062 545298 186146 545534
rect 186382 545298 221826 545534
rect 222062 545298 222146 545534
rect 222382 545298 257826 545534
rect 258062 545298 258146 545534
rect 258382 545298 293826 545534
rect 294062 545298 294146 545534
rect 294382 545298 329826 545534
rect 330062 545298 330146 545534
rect 330382 545298 365826 545534
rect 366062 545298 366146 545534
rect 366382 545298 401826 545534
rect 402062 545298 402146 545534
rect 402382 545298 570350 545534
rect 570586 545298 570670 545534
rect 570906 545298 585342 545534
rect 585578 545298 585662 545534
rect 585898 545298 592650 545534
rect -8726 545266 592650 545298
rect -8726 514354 592650 514386
rect -8726 514118 -2934 514354
rect -2698 514118 -2614 514354
rect -2378 514118 13198 514354
rect 13434 514118 13518 514354
rect 13754 514118 167826 514354
rect 168062 514118 168146 514354
rect 168382 514118 203826 514354
rect 204062 514118 204146 514354
rect 204382 514118 239826 514354
rect 240062 514118 240146 514354
rect 240382 514118 275826 514354
rect 276062 514118 276146 514354
rect 276382 514118 311826 514354
rect 312062 514118 312146 514354
rect 312382 514118 347826 514354
rect 348062 514118 348146 514354
rect 348382 514118 383826 514354
rect 384062 514118 384146 514354
rect 384382 514118 419826 514354
rect 420062 514118 420146 514354
rect 420382 514118 563826 514354
rect 564062 514118 564146 514354
rect 564382 514118 582326 514354
rect 582562 514118 582646 514354
rect 582882 514118 586302 514354
rect 586538 514118 586622 514354
rect 586858 514118 592650 514354
rect -8726 514034 592650 514118
rect -8726 513798 -2934 514034
rect -2698 513798 -2614 514034
rect -2378 513798 13198 514034
rect 13434 513798 13518 514034
rect 13754 513798 167826 514034
rect 168062 513798 168146 514034
rect 168382 513798 203826 514034
rect 204062 513798 204146 514034
rect 204382 513798 239826 514034
rect 240062 513798 240146 514034
rect 240382 513798 275826 514034
rect 276062 513798 276146 514034
rect 276382 513798 311826 514034
rect 312062 513798 312146 514034
rect 312382 513798 347826 514034
rect 348062 513798 348146 514034
rect 348382 513798 383826 514034
rect 384062 513798 384146 514034
rect 384382 513798 419826 514034
rect 420062 513798 420146 514034
rect 420382 513798 563826 514034
rect 564062 513798 564146 514034
rect 564382 513798 582326 514034
rect 582562 513798 582646 514034
rect 582882 513798 586302 514034
rect 586538 513798 586622 514034
rect 586858 513798 592650 514034
rect -8726 513766 592650 513798
rect -8726 509854 592650 509886
rect -8726 509618 -1974 509854
rect -1738 509618 -1654 509854
rect -1418 509618 5826 509854
rect 6062 509618 6146 509854
rect 6382 509618 185826 509854
rect 186062 509618 186146 509854
rect 186382 509618 221826 509854
rect 222062 509618 222146 509854
rect 222382 509618 257826 509854
rect 258062 509618 258146 509854
rect 258382 509618 293826 509854
rect 294062 509618 294146 509854
rect 294382 509618 329826 509854
rect 330062 509618 330146 509854
rect 330382 509618 365826 509854
rect 366062 509618 366146 509854
rect 366382 509618 401826 509854
rect 402062 509618 402146 509854
rect 402382 509618 570350 509854
rect 570586 509618 570670 509854
rect 570906 509618 585342 509854
rect 585578 509618 585662 509854
rect 585898 509618 592650 509854
rect -8726 509534 592650 509618
rect -8726 509298 -1974 509534
rect -1738 509298 -1654 509534
rect -1418 509298 5826 509534
rect 6062 509298 6146 509534
rect 6382 509298 185826 509534
rect 186062 509298 186146 509534
rect 186382 509298 221826 509534
rect 222062 509298 222146 509534
rect 222382 509298 257826 509534
rect 258062 509298 258146 509534
rect 258382 509298 293826 509534
rect 294062 509298 294146 509534
rect 294382 509298 329826 509534
rect 330062 509298 330146 509534
rect 330382 509298 365826 509534
rect 366062 509298 366146 509534
rect 366382 509298 401826 509534
rect 402062 509298 402146 509534
rect 402382 509298 570350 509534
rect 570586 509298 570670 509534
rect 570906 509298 585342 509534
rect 585578 509298 585662 509534
rect 585898 509298 592650 509534
rect -8726 509266 592650 509298
rect -8726 478354 592650 478386
rect -8726 478118 -2934 478354
rect -2698 478118 -2614 478354
rect -2378 478118 23826 478354
rect 24062 478118 24146 478354
rect 24382 478118 59826 478354
rect 60062 478118 60146 478354
rect 60382 478118 95826 478354
rect 96062 478118 96146 478354
rect 96382 478118 131826 478354
rect 132062 478118 132146 478354
rect 132382 478118 167826 478354
rect 168062 478118 168146 478354
rect 168382 478118 203826 478354
rect 204062 478118 204146 478354
rect 204382 478118 239826 478354
rect 240062 478118 240146 478354
rect 240382 478118 275826 478354
rect 276062 478118 276146 478354
rect 276382 478118 311826 478354
rect 312062 478118 312146 478354
rect 312382 478118 347826 478354
rect 348062 478118 348146 478354
rect 348382 478118 383826 478354
rect 384062 478118 384146 478354
rect 384382 478118 419826 478354
rect 420062 478118 420146 478354
rect 420382 478118 455826 478354
rect 456062 478118 456146 478354
rect 456382 478118 491826 478354
rect 492062 478118 492146 478354
rect 492382 478118 527826 478354
rect 528062 478118 528146 478354
rect 528382 478118 563826 478354
rect 564062 478118 564146 478354
rect 564382 478118 582326 478354
rect 582562 478118 582646 478354
rect 582882 478118 586302 478354
rect 586538 478118 586622 478354
rect 586858 478118 592650 478354
rect -8726 478034 592650 478118
rect -8726 477798 -2934 478034
rect -2698 477798 -2614 478034
rect -2378 477798 23826 478034
rect 24062 477798 24146 478034
rect 24382 477798 59826 478034
rect 60062 477798 60146 478034
rect 60382 477798 95826 478034
rect 96062 477798 96146 478034
rect 96382 477798 131826 478034
rect 132062 477798 132146 478034
rect 132382 477798 167826 478034
rect 168062 477798 168146 478034
rect 168382 477798 203826 478034
rect 204062 477798 204146 478034
rect 204382 477798 239826 478034
rect 240062 477798 240146 478034
rect 240382 477798 275826 478034
rect 276062 477798 276146 478034
rect 276382 477798 311826 478034
rect 312062 477798 312146 478034
rect 312382 477798 347826 478034
rect 348062 477798 348146 478034
rect 348382 477798 383826 478034
rect 384062 477798 384146 478034
rect 384382 477798 419826 478034
rect 420062 477798 420146 478034
rect 420382 477798 455826 478034
rect 456062 477798 456146 478034
rect 456382 477798 491826 478034
rect 492062 477798 492146 478034
rect 492382 477798 527826 478034
rect 528062 477798 528146 478034
rect 528382 477798 563826 478034
rect 564062 477798 564146 478034
rect 564382 477798 582326 478034
rect 582562 477798 582646 478034
rect 582882 477798 586302 478034
rect 586538 477798 586622 478034
rect 586858 477798 592650 478034
rect -8726 477766 592650 477798
rect -8726 473854 592650 473886
rect -8726 473618 -1974 473854
rect -1738 473618 -1654 473854
rect -1418 473618 5826 473854
rect 6062 473618 6146 473854
rect 6382 473618 41826 473854
rect 42062 473618 42146 473854
rect 42382 473618 77826 473854
rect 78062 473618 78146 473854
rect 78382 473618 113826 473854
rect 114062 473618 114146 473854
rect 114382 473618 149826 473854
rect 150062 473618 150146 473854
rect 150382 473618 185826 473854
rect 186062 473618 186146 473854
rect 186382 473618 221826 473854
rect 222062 473618 222146 473854
rect 222382 473618 257826 473854
rect 258062 473618 258146 473854
rect 258382 473618 293826 473854
rect 294062 473618 294146 473854
rect 294382 473618 329826 473854
rect 330062 473618 330146 473854
rect 330382 473618 365826 473854
rect 366062 473618 366146 473854
rect 366382 473618 401826 473854
rect 402062 473618 402146 473854
rect 402382 473618 437826 473854
rect 438062 473618 438146 473854
rect 438382 473618 473826 473854
rect 474062 473618 474146 473854
rect 474382 473618 509826 473854
rect 510062 473618 510146 473854
rect 510382 473618 545826 473854
rect 546062 473618 546146 473854
rect 546382 473618 585342 473854
rect 585578 473618 585662 473854
rect 585898 473618 592650 473854
rect -8726 473534 592650 473618
rect -8726 473298 -1974 473534
rect -1738 473298 -1654 473534
rect -1418 473298 5826 473534
rect 6062 473298 6146 473534
rect 6382 473298 41826 473534
rect 42062 473298 42146 473534
rect 42382 473298 77826 473534
rect 78062 473298 78146 473534
rect 78382 473298 113826 473534
rect 114062 473298 114146 473534
rect 114382 473298 149826 473534
rect 150062 473298 150146 473534
rect 150382 473298 185826 473534
rect 186062 473298 186146 473534
rect 186382 473298 221826 473534
rect 222062 473298 222146 473534
rect 222382 473298 257826 473534
rect 258062 473298 258146 473534
rect 258382 473298 293826 473534
rect 294062 473298 294146 473534
rect 294382 473298 329826 473534
rect 330062 473298 330146 473534
rect 330382 473298 365826 473534
rect 366062 473298 366146 473534
rect 366382 473298 401826 473534
rect 402062 473298 402146 473534
rect 402382 473298 437826 473534
rect 438062 473298 438146 473534
rect 438382 473298 473826 473534
rect 474062 473298 474146 473534
rect 474382 473298 509826 473534
rect 510062 473298 510146 473534
rect 510382 473298 545826 473534
rect 546062 473298 546146 473534
rect 546382 473298 585342 473534
rect 585578 473298 585662 473534
rect 585898 473298 592650 473534
rect -8726 473266 592650 473298
rect -8726 442354 592650 442386
rect -8726 442118 -2934 442354
rect -2698 442118 -2614 442354
rect -2378 442118 13198 442354
rect 13434 442118 13518 442354
rect 13754 442118 167826 442354
rect 168062 442118 168146 442354
rect 168382 442118 203826 442354
rect 204062 442118 204146 442354
rect 204382 442118 239826 442354
rect 240062 442118 240146 442354
rect 240382 442118 275826 442354
rect 276062 442118 276146 442354
rect 276382 442118 311826 442354
rect 312062 442118 312146 442354
rect 312382 442118 347826 442354
rect 348062 442118 348146 442354
rect 348382 442118 383826 442354
rect 384062 442118 384146 442354
rect 384382 442118 419826 442354
rect 420062 442118 420146 442354
rect 420382 442118 563826 442354
rect 564062 442118 564146 442354
rect 564382 442118 582326 442354
rect 582562 442118 582646 442354
rect 582882 442118 586302 442354
rect 586538 442118 586622 442354
rect 586858 442118 592650 442354
rect -8726 442034 592650 442118
rect -8726 441798 -2934 442034
rect -2698 441798 -2614 442034
rect -2378 441798 13198 442034
rect 13434 441798 13518 442034
rect 13754 441798 167826 442034
rect 168062 441798 168146 442034
rect 168382 441798 203826 442034
rect 204062 441798 204146 442034
rect 204382 441798 239826 442034
rect 240062 441798 240146 442034
rect 240382 441798 275826 442034
rect 276062 441798 276146 442034
rect 276382 441798 311826 442034
rect 312062 441798 312146 442034
rect 312382 441798 347826 442034
rect 348062 441798 348146 442034
rect 348382 441798 383826 442034
rect 384062 441798 384146 442034
rect 384382 441798 419826 442034
rect 420062 441798 420146 442034
rect 420382 441798 563826 442034
rect 564062 441798 564146 442034
rect 564382 441798 582326 442034
rect 582562 441798 582646 442034
rect 582882 441798 586302 442034
rect 586538 441798 586622 442034
rect 586858 441798 592650 442034
rect -8726 441766 592650 441798
rect -8726 437854 592650 437886
rect -8726 437618 -1974 437854
rect -1738 437618 -1654 437854
rect -1418 437618 5826 437854
rect 6062 437618 6146 437854
rect 6382 437618 185826 437854
rect 186062 437618 186146 437854
rect 186382 437618 221826 437854
rect 222062 437618 222146 437854
rect 222382 437618 257826 437854
rect 258062 437618 258146 437854
rect 258382 437618 293826 437854
rect 294062 437618 294146 437854
rect 294382 437618 329826 437854
rect 330062 437618 330146 437854
rect 330382 437618 365826 437854
rect 366062 437618 366146 437854
rect 366382 437618 401826 437854
rect 402062 437618 402146 437854
rect 402382 437618 570350 437854
rect 570586 437618 570670 437854
rect 570906 437618 585342 437854
rect 585578 437618 585662 437854
rect 585898 437618 592650 437854
rect -8726 437534 592650 437618
rect -8726 437298 -1974 437534
rect -1738 437298 -1654 437534
rect -1418 437298 5826 437534
rect 6062 437298 6146 437534
rect 6382 437298 185826 437534
rect 186062 437298 186146 437534
rect 186382 437298 221826 437534
rect 222062 437298 222146 437534
rect 222382 437298 257826 437534
rect 258062 437298 258146 437534
rect 258382 437298 293826 437534
rect 294062 437298 294146 437534
rect 294382 437298 329826 437534
rect 330062 437298 330146 437534
rect 330382 437298 365826 437534
rect 366062 437298 366146 437534
rect 366382 437298 401826 437534
rect 402062 437298 402146 437534
rect 402382 437298 570350 437534
rect 570586 437298 570670 437534
rect 570906 437298 585342 437534
rect 585578 437298 585662 437534
rect 585898 437298 592650 437534
rect -8726 437266 592650 437298
rect -8726 406354 592650 406386
rect -8726 406118 -2934 406354
rect -2698 406118 -2614 406354
rect -2378 406118 13198 406354
rect 13434 406118 13518 406354
rect 13754 406118 167826 406354
rect 168062 406118 168146 406354
rect 168382 406118 203826 406354
rect 204062 406118 204146 406354
rect 204382 406118 239826 406354
rect 240062 406118 240146 406354
rect 240382 406118 275826 406354
rect 276062 406118 276146 406354
rect 276382 406118 311826 406354
rect 312062 406118 312146 406354
rect 312382 406118 347826 406354
rect 348062 406118 348146 406354
rect 348382 406118 383826 406354
rect 384062 406118 384146 406354
rect 384382 406118 419826 406354
rect 420062 406118 420146 406354
rect 420382 406118 563826 406354
rect 564062 406118 564146 406354
rect 564382 406118 582326 406354
rect 582562 406118 582646 406354
rect 582882 406118 586302 406354
rect 586538 406118 586622 406354
rect 586858 406118 592650 406354
rect -8726 406034 592650 406118
rect -8726 405798 -2934 406034
rect -2698 405798 -2614 406034
rect -2378 405798 13198 406034
rect 13434 405798 13518 406034
rect 13754 405798 167826 406034
rect 168062 405798 168146 406034
rect 168382 405798 203826 406034
rect 204062 405798 204146 406034
rect 204382 405798 239826 406034
rect 240062 405798 240146 406034
rect 240382 405798 275826 406034
rect 276062 405798 276146 406034
rect 276382 405798 311826 406034
rect 312062 405798 312146 406034
rect 312382 405798 347826 406034
rect 348062 405798 348146 406034
rect 348382 405798 383826 406034
rect 384062 405798 384146 406034
rect 384382 405798 419826 406034
rect 420062 405798 420146 406034
rect 420382 405798 563826 406034
rect 564062 405798 564146 406034
rect 564382 405798 582326 406034
rect 582562 405798 582646 406034
rect 582882 405798 586302 406034
rect 586538 405798 586622 406034
rect 586858 405798 592650 406034
rect -8726 405766 592650 405798
rect -8726 401854 592650 401886
rect -8726 401618 -1974 401854
rect -1738 401618 -1654 401854
rect -1418 401618 5826 401854
rect 6062 401618 6146 401854
rect 6382 401618 185826 401854
rect 186062 401618 186146 401854
rect 186382 401618 221826 401854
rect 222062 401618 222146 401854
rect 222382 401618 257826 401854
rect 258062 401618 258146 401854
rect 258382 401618 293826 401854
rect 294062 401618 294146 401854
rect 294382 401618 329826 401854
rect 330062 401618 330146 401854
rect 330382 401618 365826 401854
rect 366062 401618 366146 401854
rect 366382 401618 401826 401854
rect 402062 401618 402146 401854
rect 402382 401618 570350 401854
rect 570586 401618 570670 401854
rect 570906 401618 585342 401854
rect 585578 401618 585662 401854
rect 585898 401618 592650 401854
rect -8726 401534 592650 401618
rect -8726 401298 -1974 401534
rect -1738 401298 -1654 401534
rect -1418 401298 5826 401534
rect 6062 401298 6146 401534
rect 6382 401298 185826 401534
rect 186062 401298 186146 401534
rect 186382 401298 221826 401534
rect 222062 401298 222146 401534
rect 222382 401298 257826 401534
rect 258062 401298 258146 401534
rect 258382 401298 293826 401534
rect 294062 401298 294146 401534
rect 294382 401298 329826 401534
rect 330062 401298 330146 401534
rect 330382 401298 365826 401534
rect 366062 401298 366146 401534
rect 366382 401298 401826 401534
rect 402062 401298 402146 401534
rect 402382 401298 570350 401534
rect 570586 401298 570670 401534
rect 570906 401298 585342 401534
rect 585578 401298 585662 401534
rect 585898 401298 592650 401534
rect -8726 401266 592650 401298
rect -8726 370354 592650 370386
rect -8726 370118 -2934 370354
rect -2698 370118 -2614 370354
rect -2378 370118 13198 370354
rect 13434 370118 13518 370354
rect 13754 370118 167826 370354
rect 168062 370118 168146 370354
rect 168382 370118 203826 370354
rect 204062 370118 204146 370354
rect 204382 370118 239826 370354
rect 240062 370118 240146 370354
rect 240382 370118 275826 370354
rect 276062 370118 276146 370354
rect 276382 370118 311826 370354
rect 312062 370118 312146 370354
rect 312382 370118 347826 370354
rect 348062 370118 348146 370354
rect 348382 370118 383826 370354
rect 384062 370118 384146 370354
rect 384382 370118 419826 370354
rect 420062 370118 420146 370354
rect 420382 370118 563826 370354
rect 564062 370118 564146 370354
rect 564382 370118 582326 370354
rect 582562 370118 582646 370354
rect 582882 370118 586302 370354
rect 586538 370118 586622 370354
rect 586858 370118 592650 370354
rect -8726 370034 592650 370118
rect -8726 369798 -2934 370034
rect -2698 369798 -2614 370034
rect -2378 369798 13198 370034
rect 13434 369798 13518 370034
rect 13754 369798 167826 370034
rect 168062 369798 168146 370034
rect 168382 369798 203826 370034
rect 204062 369798 204146 370034
rect 204382 369798 239826 370034
rect 240062 369798 240146 370034
rect 240382 369798 275826 370034
rect 276062 369798 276146 370034
rect 276382 369798 311826 370034
rect 312062 369798 312146 370034
rect 312382 369798 347826 370034
rect 348062 369798 348146 370034
rect 348382 369798 383826 370034
rect 384062 369798 384146 370034
rect 384382 369798 419826 370034
rect 420062 369798 420146 370034
rect 420382 369798 563826 370034
rect 564062 369798 564146 370034
rect 564382 369798 582326 370034
rect 582562 369798 582646 370034
rect 582882 369798 586302 370034
rect 586538 369798 586622 370034
rect 586858 369798 592650 370034
rect -8726 369766 592650 369798
rect -8726 365854 592650 365886
rect -8726 365618 -1974 365854
rect -1738 365618 -1654 365854
rect -1418 365618 5826 365854
rect 6062 365618 6146 365854
rect 6382 365618 41826 365854
rect 42062 365618 42146 365854
rect 42382 365618 77826 365854
rect 78062 365618 78146 365854
rect 78382 365618 113826 365854
rect 114062 365618 114146 365854
rect 114382 365618 149826 365854
rect 150062 365618 150146 365854
rect 150382 365618 185826 365854
rect 186062 365618 186146 365854
rect 186382 365618 221826 365854
rect 222062 365618 222146 365854
rect 222382 365618 257826 365854
rect 258062 365618 258146 365854
rect 258382 365618 293826 365854
rect 294062 365618 294146 365854
rect 294382 365618 329826 365854
rect 330062 365618 330146 365854
rect 330382 365618 365826 365854
rect 366062 365618 366146 365854
rect 366382 365618 401826 365854
rect 402062 365618 402146 365854
rect 402382 365618 437826 365854
rect 438062 365618 438146 365854
rect 438382 365618 473826 365854
rect 474062 365618 474146 365854
rect 474382 365618 509826 365854
rect 510062 365618 510146 365854
rect 510382 365618 545826 365854
rect 546062 365618 546146 365854
rect 546382 365618 585342 365854
rect 585578 365618 585662 365854
rect 585898 365618 592650 365854
rect -8726 365534 592650 365618
rect -8726 365298 -1974 365534
rect -1738 365298 -1654 365534
rect -1418 365298 5826 365534
rect 6062 365298 6146 365534
rect 6382 365298 41826 365534
rect 42062 365298 42146 365534
rect 42382 365298 77826 365534
rect 78062 365298 78146 365534
rect 78382 365298 113826 365534
rect 114062 365298 114146 365534
rect 114382 365298 149826 365534
rect 150062 365298 150146 365534
rect 150382 365298 185826 365534
rect 186062 365298 186146 365534
rect 186382 365298 221826 365534
rect 222062 365298 222146 365534
rect 222382 365298 257826 365534
rect 258062 365298 258146 365534
rect 258382 365298 293826 365534
rect 294062 365298 294146 365534
rect 294382 365298 329826 365534
rect 330062 365298 330146 365534
rect 330382 365298 365826 365534
rect 366062 365298 366146 365534
rect 366382 365298 401826 365534
rect 402062 365298 402146 365534
rect 402382 365298 437826 365534
rect 438062 365298 438146 365534
rect 438382 365298 473826 365534
rect 474062 365298 474146 365534
rect 474382 365298 509826 365534
rect 510062 365298 510146 365534
rect 510382 365298 545826 365534
rect 546062 365298 546146 365534
rect 546382 365298 585342 365534
rect 585578 365298 585662 365534
rect 585898 365298 592650 365534
rect -8726 365266 592650 365298
rect -8726 334354 592650 334386
rect -8726 334118 -2934 334354
rect -2698 334118 -2614 334354
rect -2378 334118 13198 334354
rect 13434 334118 13518 334354
rect 13754 334118 167826 334354
rect 168062 334118 168146 334354
rect 168382 334118 203826 334354
rect 204062 334118 204146 334354
rect 204382 334118 239826 334354
rect 240062 334118 240146 334354
rect 240382 334118 275826 334354
rect 276062 334118 276146 334354
rect 276382 334118 311826 334354
rect 312062 334118 312146 334354
rect 312382 334118 347826 334354
rect 348062 334118 348146 334354
rect 348382 334118 383826 334354
rect 384062 334118 384146 334354
rect 384382 334118 419826 334354
rect 420062 334118 420146 334354
rect 420382 334118 563826 334354
rect 564062 334118 564146 334354
rect 564382 334118 582326 334354
rect 582562 334118 582646 334354
rect 582882 334118 586302 334354
rect 586538 334118 586622 334354
rect 586858 334118 592650 334354
rect -8726 334034 592650 334118
rect -8726 333798 -2934 334034
rect -2698 333798 -2614 334034
rect -2378 333798 13198 334034
rect 13434 333798 13518 334034
rect 13754 333798 167826 334034
rect 168062 333798 168146 334034
rect 168382 333798 203826 334034
rect 204062 333798 204146 334034
rect 204382 333798 239826 334034
rect 240062 333798 240146 334034
rect 240382 333798 275826 334034
rect 276062 333798 276146 334034
rect 276382 333798 311826 334034
rect 312062 333798 312146 334034
rect 312382 333798 347826 334034
rect 348062 333798 348146 334034
rect 348382 333798 383826 334034
rect 384062 333798 384146 334034
rect 384382 333798 419826 334034
rect 420062 333798 420146 334034
rect 420382 333798 563826 334034
rect 564062 333798 564146 334034
rect 564382 333798 582326 334034
rect 582562 333798 582646 334034
rect 582882 333798 586302 334034
rect 586538 333798 586622 334034
rect 586858 333798 592650 334034
rect -8726 333766 592650 333798
rect -8726 329854 592650 329886
rect -8726 329618 -1974 329854
rect -1738 329618 -1654 329854
rect -1418 329618 5826 329854
rect 6062 329618 6146 329854
rect 6382 329618 185826 329854
rect 186062 329618 186146 329854
rect 186382 329618 221826 329854
rect 222062 329618 222146 329854
rect 222382 329618 257826 329854
rect 258062 329618 258146 329854
rect 258382 329618 293826 329854
rect 294062 329618 294146 329854
rect 294382 329618 329826 329854
rect 330062 329618 330146 329854
rect 330382 329618 365826 329854
rect 366062 329618 366146 329854
rect 366382 329618 401826 329854
rect 402062 329618 402146 329854
rect 402382 329618 570350 329854
rect 570586 329618 570670 329854
rect 570906 329618 585342 329854
rect 585578 329618 585662 329854
rect 585898 329618 592650 329854
rect -8726 329534 592650 329618
rect -8726 329298 -1974 329534
rect -1738 329298 -1654 329534
rect -1418 329298 5826 329534
rect 6062 329298 6146 329534
rect 6382 329298 185826 329534
rect 186062 329298 186146 329534
rect 186382 329298 221826 329534
rect 222062 329298 222146 329534
rect 222382 329298 257826 329534
rect 258062 329298 258146 329534
rect 258382 329298 293826 329534
rect 294062 329298 294146 329534
rect 294382 329298 329826 329534
rect 330062 329298 330146 329534
rect 330382 329298 365826 329534
rect 366062 329298 366146 329534
rect 366382 329298 401826 329534
rect 402062 329298 402146 329534
rect 402382 329298 570350 329534
rect 570586 329298 570670 329534
rect 570906 329298 585342 329534
rect 585578 329298 585662 329534
rect 585898 329298 592650 329534
rect -8726 329266 592650 329298
rect -8726 298354 592650 298386
rect -8726 298118 -2934 298354
rect -2698 298118 -2614 298354
rect -2378 298118 13198 298354
rect 13434 298118 13518 298354
rect 13754 298118 167826 298354
rect 168062 298118 168146 298354
rect 168382 298118 203826 298354
rect 204062 298118 204146 298354
rect 204382 298118 239826 298354
rect 240062 298118 240146 298354
rect 240382 298118 275826 298354
rect 276062 298118 276146 298354
rect 276382 298118 311826 298354
rect 312062 298118 312146 298354
rect 312382 298118 347826 298354
rect 348062 298118 348146 298354
rect 348382 298118 383826 298354
rect 384062 298118 384146 298354
rect 384382 298118 419826 298354
rect 420062 298118 420146 298354
rect 420382 298118 563826 298354
rect 564062 298118 564146 298354
rect 564382 298118 582326 298354
rect 582562 298118 582646 298354
rect 582882 298118 586302 298354
rect 586538 298118 586622 298354
rect 586858 298118 592650 298354
rect -8726 298034 592650 298118
rect -8726 297798 -2934 298034
rect -2698 297798 -2614 298034
rect -2378 297798 13198 298034
rect 13434 297798 13518 298034
rect 13754 297798 167826 298034
rect 168062 297798 168146 298034
rect 168382 297798 203826 298034
rect 204062 297798 204146 298034
rect 204382 297798 239826 298034
rect 240062 297798 240146 298034
rect 240382 297798 275826 298034
rect 276062 297798 276146 298034
rect 276382 297798 311826 298034
rect 312062 297798 312146 298034
rect 312382 297798 347826 298034
rect 348062 297798 348146 298034
rect 348382 297798 383826 298034
rect 384062 297798 384146 298034
rect 384382 297798 419826 298034
rect 420062 297798 420146 298034
rect 420382 297798 563826 298034
rect 564062 297798 564146 298034
rect 564382 297798 582326 298034
rect 582562 297798 582646 298034
rect 582882 297798 586302 298034
rect 586538 297798 586622 298034
rect 586858 297798 592650 298034
rect -8726 297766 592650 297798
rect -8726 293854 592650 293886
rect -8726 293618 -1974 293854
rect -1738 293618 -1654 293854
rect -1418 293618 5826 293854
rect 6062 293618 6146 293854
rect 6382 293618 185826 293854
rect 186062 293618 186146 293854
rect 186382 293618 221826 293854
rect 222062 293618 222146 293854
rect 222382 293618 257826 293854
rect 258062 293618 258146 293854
rect 258382 293618 293826 293854
rect 294062 293618 294146 293854
rect 294382 293618 329826 293854
rect 330062 293618 330146 293854
rect 330382 293618 365826 293854
rect 366062 293618 366146 293854
rect 366382 293618 401826 293854
rect 402062 293618 402146 293854
rect 402382 293618 570350 293854
rect 570586 293618 570670 293854
rect 570906 293618 585342 293854
rect 585578 293618 585662 293854
rect 585898 293618 592650 293854
rect -8726 293534 592650 293618
rect -8726 293298 -1974 293534
rect -1738 293298 -1654 293534
rect -1418 293298 5826 293534
rect 6062 293298 6146 293534
rect 6382 293298 185826 293534
rect 186062 293298 186146 293534
rect 186382 293298 221826 293534
rect 222062 293298 222146 293534
rect 222382 293298 257826 293534
rect 258062 293298 258146 293534
rect 258382 293298 293826 293534
rect 294062 293298 294146 293534
rect 294382 293298 329826 293534
rect 330062 293298 330146 293534
rect 330382 293298 365826 293534
rect 366062 293298 366146 293534
rect 366382 293298 401826 293534
rect 402062 293298 402146 293534
rect 402382 293298 570350 293534
rect 570586 293298 570670 293534
rect 570906 293298 585342 293534
rect 585578 293298 585662 293534
rect 585898 293298 592650 293534
rect -8726 293266 592650 293298
rect -8726 262354 592650 262386
rect -8726 262118 -2934 262354
rect -2698 262118 -2614 262354
rect -2378 262118 13198 262354
rect 13434 262118 13518 262354
rect 13754 262118 167826 262354
rect 168062 262118 168146 262354
rect 168382 262118 203826 262354
rect 204062 262118 204146 262354
rect 204382 262118 239826 262354
rect 240062 262118 240146 262354
rect 240382 262118 275826 262354
rect 276062 262118 276146 262354
rect 276382 262118 311826 262354
rect 312062 262118 312146 262354
rect 312382 262118 347826 262354
rect 348062 262118 348146 262354
rect 348382 262118 383826 262354
rect 384062 262118 384146 262354
rect 384382 262118 419826 262354
rect 420062 262118 420146 262354
rect 420382 262118 563826 262354
rect 564062 262118 564146 262354
rect 564382 262118 582326 262354
rect 582562 262118 582646 262354
rect 582882 262118 586302 262354
rect 586538 262118 586622 262354
rect 586858 262118 592650 262354
rect -8726 262034 592650 262118
rect -8726 261798 -2934 262034
rect -2698 261798 -2614 262034
rect -2378 261798 13198 262034
rect 13434 261798 13518 262034
rect 13754 261798 167826 262034
rect 168062 261798 168146 262034
rect 168382 261798 203826 262034
rect 204062 261798 204146 262034
rect 204382 261798 239826 262034
rect 240062 261798 240146 262034
rect 240382 261798 275826 262034
rect 276062 261798 276146 262034
rect 276382 261798 311826 262034
rect 312062 261798 312146 262034
rect 312382 261798 347826 262034
rect 348062 261798 348146 262034
rect 348382 261798 383826 262034
rect 384062 261798 384146 262034
rect 384382 261798 419826 262034
rect 420062 261798 420146 262034
rect 420382 261798 563826 262034
rect 564062 261798 564146 262034
rect 564382 261798 582326 262034
rect 582562 261798 582646 262034
rect 582882 261798 586302 262034
rect 586538 261798 586622 262034
rect 586858 261798 592650 262034
rect -8726 261766 592650 261798
rect -8726 257854 592650 257886
rect -8726 257618 -1974 257854
rect -1738 257618 -1654 257854
rect -1418 257618 5826 257854
rect 6062 257618 6146 257854
rect 6382 257618 185826 257854
rect 186062 257618 186146 257854
rect 186382 257618 221826 257854
rect 222062 257618 222146 257854
rect 222382 257618 257826 257854
rect 258062 257618 258146 257854
rect 258382 257618 293826 257854
rect 294062 257618 294146 257854
rect 294382 257618 329826 257854
rect 330062 257618 330146 257854
rect 330382 257618 365826 257854
rect 366062 257618 366146 257854
rect 366382 257618 401826 257854
rect 402062 257618 402146 257854
rect 402382 257618 570350 257854
rect 570586 257618 570670 257854
rect 570906 257618 585342 257854
rect 585578 257618 585662 257854
rect 585898 257618 592650 257854
rect -8726 257534 592650 257618
rect -8726 257298 -1974 257534
rect -1738 257298 -1654 257534
rect -1418 257298 5826 257534
rect 6062 257298 6146 257534
rect 6382 257298 185826 257534
rect 186062 257298 186146 257534
rect 186382 257298 221826 257534
rect 222062 257298 222146 257534
rect 222382 257298 257826 257534
rect 258062 257298 258146 257534
rect 258382 257298 293826 257534
rect 294062 257298 294146 257534
rect 294382 257298 329826 257534
rect 330062 257298 330146 257534
rect 330382 257298 365826 257534
rect 366062 257298 366146 257534
rect 366382 257298 401826 257534
rect 402062 257298 402146 257534
rect 402382 257298 570350 257534
rect 570586 257298 570670 257534
rect 570906 257298 585342 257534
rect 585578 257298 585662 257534
rect 585898 257298 592650 257534
rect -8726 257266 592650 257298
rect -8726 226354 592650 226386
rect -8726 226118 -2934 226354
rect -2698 226118 -2614 226354
rect -2378 226118 13198 226354
rect 13434 226118 13518 226354
rect 13754 226118 167826 226354
rect 168062 226118 168146 226354
rect 168382 226118 203826 226354
rect 204062 226118 204146 226354
rect 204382 226118 239826 226354
rect 240062 226118 240146 226354
rect 240382 226118 275826 226354
rect 276062 226118 276146 226354
rect 276382 226118 311826 226354
rect 312062 226118 312146 226354
rect 312382 226118 347826 226354
rect 348062 226118 348146 226354
rect 348382 226118 383826 226354
rect 384062 226118 384146 226354
rect 384382 226118 419826 226354
rect 420062 226118 420146 226354
rect 420382 226118 563826 226354
rect 564062 226118 564146 226354
rect 564382 226118 582326 226354
rect 582562 226118 582646 226354
rect 582882 226118 586302 226354
rect 586538 226118 586622 226354
rect 586858 226118 592650 226354
rect -8726 226034 592650 226118
rect -8726 225798 -2934 226034
rect -2698 225798 -2614 226034
rect -2378 225798 13198 226034
rect 13434 225798 13518 226034
rect 13754 225798 167826 226034
rect 168062 225798 168146 226034
rect 168382 225798 203826 226034
rect 204062 225798 204146 226034
rect 204382 225798 239826 226034
rect 240062 225798 240146 226034
rect 240382 225798 275826 226034
rect 276062 225798 276146 226034
rect 276382 225798 311826 226034
rect 312062 225798 312146 226034
rect 312382 225798 347826 226034
rect 348062 225798 348146 226034
rect 348382 225798 383826 226034
rect 384062 225798 384146 226034
rect 384382 225798 419826 226034
rect 420062 225798 420146 226034
rect 420382 225798 563826 226034
rect 564062 225798 564146 226034
rect 564382 225798 582326 226034
rect 582562 225798 582646 226034
rect 582882 225798 586302 226034
rect 586538 225798 586622 226034
rect 586858 225798 592650 226034
rect -8726 225766 592650 225798
rect -8726 221854 592650 221886
rect -8726 221618 -1974 221854
rect -1738 221618 -1654 221854
rect -1418 221618 5826 221854
rect 6062 221618 6146 221854
rect 6382 221618 185826 221854
rect 186062 221618 186146 221854
rect 186382 221618 221826 221854
rect 222062 221618 222146 221854
rect 222382 221618 257826 221854
rect 258062 221618 258146 221854
rect 258382 221618 293826 221854
rect 294062 221618 294146 221854
rect 294382 221618 329826 221854
rect 330062 221618 330146 221854
rect 330382 221618 365826 221854
rect 366062 221618 366146 221854
rect 366382 221618 401826 221854
rect 402062 221618 402146 221854
rect 402382 221618 570350 221854
rect 570586 221618 570670 221854
rect 570906 221618 585342 221854
rect 585578 221618 585662 221854
rect 585898 221618 592650 221854
rect -8726 221534 592650 221618
rect -8726 221298 -1974 221534
rect -1738 221298 -1654 221534
rect -1418 221298 5826 221534
rect 6062 221298 6146 221534
rect 6382 221298 185826 221534
rect 186062 221298 186146 221534
rect 186382 221298 221826 221534
rect 222062 221298 222146 221534
rect 222382 221298 257826 221534
rect 258062 221298 258146 221534
rect 258382 221298 293826 221534
rect 294062 221298 294146 221534
rect 294382 221298 329826 221534
rect 330062 221298 330146 221534
rect 330382 221298 365826 221534
rect 366062 221298 366146 221534
rect 366382 221298 401826 221534
rect 402062 221298 402146 221534
rect 402382 221298 570350 221534
rect 570586 221298 570670 221534
rect 570906 221298 585342 221534
rect 585578 221298 585662 221534
rect 585898 221298 592650 221534
rect -8726 221266 592650 221298
rect -8726 190354 592650 190386
rect -8726 190118 -2934 190354
rect -2698 190118 -2614 190354
rect -2378 190118 13198 190354
rect 13434 190118 13518 190354
rect 13754 190118 167826 190354
rect 168062 190118 168146 190354
rect 168382 190118 203826 190354
rect 204062 190118 204146 190354
rect 204382 190118 239826 190354
rect 240062 190118 240146 190354
rect 240382 190118 275826 190354
rect 276062 190118 276146 190354
rect 276382 190118 311826 190354
rect 312062 190118 312146 190354
rect 312382 190118 347826 190354
rect 348062 190118 348146 190354
rect 348382 190118 383826 190354
rect 384062 190118 384146 190354
rect 384382 190118 419826 190354
rect 420062 190118 420146 190354
rect 420382 190118 563826 190354
rect 564062 190118 564146 190354
rect 564382 190118 582326 190354
rect 582562 190118 582646 190354
rect 582882 190118 586302 190354
rect 586538 190118 586622 190354
rect 586858 190118 592650 190354
rect -8726 190034 592650 190118
rect -8726 189798 -2934 190034
rect -2698 189798 -2614 190034
rect -2378 189798 13198 190034
rect 13434 189798 13518 190034
rect 13754 189798 167826 190034
rect 168062 189798 168146 190034
rect 168382 189798 203826 190034
rect 204062 189798 204146 190034
rect 204382 189798 239826 190034
rect 240062 189798 240146 190034
rect 240382 189798 275826 190034
rect 276062 189798 276146 190034
rect 276382 189798 311826 190034
rect 312062 189798 312146 190034
rect 312382 189798 347826 190034
rect 348062 189798 348146 190034
rect 348382 189798 383826 190034
rect 384062 189798 384146 190034
rect 384382 189798 419826 190034
rect 420062 189798 420146 190034
rect 420382 189798 563826 190034
rect 564062 189798 564146 190034
rect 564382 189798 582326 190034
rect 582562 189798 582646 190034
rect 582882 189798 586302 190034
rect 586538 189798 586622 190034
rect 586858 189798 592650 190034
rect -8726 189766 592650 189798
rect -8726 185854 592650 185886
rect -8726 185618 -1974 185854
rect -1738 185618 -1654 185854
rect -1418 185618 5826 185854
rect 6062 185618 6146 185854
rect 6382 185618 185826 185854
rect 186062 185618 186146 185854
rect 186382 185618 221826 185854
rect 222062 185618 222146 185854
rect 222382 185618 257826 185854
rect 258062 185618 258146 185854
rect 258382 185618 293826 185854
rect 294062 185618 294146 185854
rect 294382 185618 329826 185854
rect 330062 185618 330146 185854
rect 330382 185618 365826 185854
rect 366062 185618 366146 185854
rect 366382 185618 401826 185854
rect 402062 185618 402146 185854
rect 402382 185618 570350 185854
rect 570586 185618 570670 185854
rect 570906 185618 585342 185854
rect 585578 185618 585662 185854
rect 585898 185618 592650 185854
rect -8726 185534 592650 185618
rect -8726 185298 -1974 185534
rect -1738 185298 -1654 185534
rect -1418 185298 5826 185534
rect 6062 185298 6146 185534
rect 6382 185298 185826 185534
rect 186062 185298 186146 185534
rect 186382 185298 221826 185534
rect 222062 185298 222146 185534
rect 222382 185298 257826 185534
rect 258062 185298 258146 185534
rect 258382 185298 293826 185534
rect 294062 185298 294146 185534
rect 294382 185298 329826 185534
rect 330062 185298 330146 185534
rect 330382 185298 365826 185534
rect 366062 185298 366146 185534
rect 366382 185298 401826 185534
rect 402062 185298 402146 185534
rect 402382 185298 570350 185534
rect 570586 185298 570670 185534
rect 570906 185298 585342 185534
rect 585578 185298 585662 185534
rect 585898 185298 592650 185534
rect -8726 185266 592650 185298
rect -8726 154354 592650 154386
rect -8726 154118 -2934 154354
rect -2698 154118 -2614 154354
rect -2378 154118 13198 154354
rect 13434 154118 13518 154354
rect 13754 154118 167826 154354
rect 168062 154118 168146 154354
rect 168382 154118 203826 154354
rect 204062 154118 204146 154354
rect 204382 154118 239826 154354
rect 240062 154118 240146 154354
rect 240382 154118 275826 154354
rect 276062 154118 276146 154354
rect 276382 154118 311826 154354
rect 312062 154118 312146 154354
rect 312382 154118 347826 154354
rect 348062 154118 348146 154354
rect 348382 154118 383826 154354
rect 384062 154118 384146 154354
rect 384382 154118 419826 154354
rect 420062 154118 420146 154354
rect 420382 154118 563826 154354
rect 564062 154118 564146 154354
rect 564382 154118 582326 154354
rect 582562 154118 582646 154354
rect 582882 154118 586302 154354
rect 586538 154118 586622 154354
rect 586858 154118 592650 154354
rect -8726 154034 592650 154118
rect -8726 153798 -2934 154034
rect -2698 153798 -2614 154034
rect -2378 153798 13198 154034
rect 13434 153798 13518 154034
rect 13754 153798 167826 154034
rect 168062 153798 168146 154034
rect 168382 153798 203826 154034
rect 204062 153798 204146 154034
rect 204382 153798 239826 154034
rect 240062 153798 240146 154034
rect 240382 153798 275826 154034
rect 276062 153798 276146 154034
rect 276382 153798 311826 154034
rect 312062 153798 312146 154034
rect 312382 153798 347826 154034
rect 348062 153798 348146 154034
rect 348382 153798 383826 154034
rect 384062 153798 384146 154034
rect 384382 153798 419826 154034
rect 420062 153798 420146 154034
rect 420382 153798 563826 154034
rect 564062 153798 564146 154034
rect 564382 153798 582326 154034
rect 582562 153798 582646 154034
rect 582882 153798 586302 154034
rect 586538 153798 586622 154034
rect 586858 153798 592650 154034
rect -8726 153766 592650 153798
rect -8726 149854 592650 149886
rect -8726 149618 -1974 149854
rect -1738 149618 -1654 149854
rect -1418 149618 5826 149854
rect 6062 149618 6146 149854
rect 6382 149618 185826 149854
rect 186062 149618 186146 149854
rect 186382 149618 221826 149854
rect 222062 149618 222146 149854
rect 222382 149618 257826 149854
rect 258062 149618 258146 149854
rect 258382 149618 293826 149854
rect 294062 149618 294146 149854
rect 294382 149618 329826 149854
rect 330062 149618 330146 149854
rect 330382 149618 365826 149854
rect 366062 149618 366146 149854
rect 366382 149618 401826 149854
rect 402062 149618 402146 149854
rect 402382 149618 570350 149854
rect 570586 149618 570670 149854
rect 570906 149618 585342 149854
rect 585578 149618 585662 149854
rect 585898 149618 592650 149854
rect -8726 149534 592650 149618
rect -8726 149298 -1974 149534
rect -1738 149298 -1654 149534
rect -1418 149298 5826 149534
rect 6062 149298 6146 149534
rect 6382 149298 185826 149534
rect 186062 149298 186146 149534
rect 186382 149298 221826 149534
rect 222062 149298 222146 149534
rect 222382 149298 257826 149534
rect 258062 149298 258146 149534
rect 258382 149298 293826 149534
rect 294062 149298 294146 149534
rect 294382 149298 329826 149534
rect 330062 149298 330146 149534
rect 330382 149298 365826 149534
rect 366062 149298 366146 149534
rect 366382 149298 401826 149534
rect 402062 149298 402146 149534
rect 402382 149298 570350 149534
rect 570586 149298 570670 149534
rect 570906 149298 585342 149534
rect 585578 149298 585662 149534
rect 585898 149298 592650 149534
rect -8726 149266 592650 149298
rect -8726 118354 592650 118386
rect -8726 118118 -2934 118354
rect -2698 118118 -2614 118354
rect -2378 118118 13198 118354
rect 13434 118118 13518 118354
rect 13754 118118 167826 118354
rect 168062 118118 168146 118354
rect 168382 118118 203826 118354
rect 204062 118118 204146 118354
rect 204382 118118 239826 118354
rect 240062 118118 240146 118354
rect 240382 118118 275826 118354
rect 276062 118118 276146 118354
rect 276382 118118 311826 118354
rect 312062 118118 312146 118354
rect 312382 118118 347826 118354
rect 348062 118118 348146 118354
rect 348382 118118 383826 118354
rect 384062 118118 384146 118354
rect 384382 118118 419826 118354
rect 420062 118118 420146 118354
rect 420382 118118 563826 118354
rect 564062 118118 564146 118354
rect 564382 118118 582326 118354
rect 582562 118118 582646 118354
rect 582882 118118 586302 118354
rect 586538 118118 586622 118354
rect 586858 118118 592650 118354
rect -8726 118034 592650 118118
rect -8726 117798 -2934 118034
rect -2698 117798 -2614 118034
rect -2378 117798 13198 118034
rect 13434 117798 13518 118034
rect 13754 117798 167826 118034
rect 168062 117798 168146 118034
rect 168382 117798 203826 118034
rect 204062 117798 204146 118034
rect 204382 117798 239826 118034
rect 240062 117798 240146 118034
rect 240382 117798 275826 118034
rect 276062 117798 276146 118034
rect 276382 117798 311826 118034
rect 312062 117798 312146 118034
rect 312382 117798 347826 118034
rect 348062 117798 348146 118034
rect 348382 117798 383826 118034
rect 384062 117798 384146 118034
rect 384382 117798 419826 118034
rect 420062 117798 420146 118034
rect 420382 117798 563826 118034
rect 564062 117798 564146 118034
rect 564382 117798 582326 118034
rect 582562 117798 582646 118034
rect 582882 117798 586302 118034
rect 586538 117798 586622 118034
rect 586858 117798 592650 118034
rect -8726 117766 592650 117798
rect -8726 113854 592650 113886
rect -8726 113618 -1974 113854
rect -1738 113618 -1654 113854
rect -1418 113618 5826 113854
rect 6062 113618 6146 113854
rect 6382 113618 173094 113854
rect 173330 113618 173414 113854
rect 173650 113618 293826 113854
rect 294062 113618 294146 113854
rect 294382 113618 401826 113854
rect 402062 113618 402146 113854
rect 402382 113618 570350 113854
rect 570586 113618 570670 113854
rect 570906 113618 585342 113854
rect 585578 113618 585662 113854
rect 585898 113618 592650 113854
rect -8726 113534 592650 113618
rect -8726 113298 -1974 113534
rect -1738 113298 -1654 113534
rect -1418 113298 5826 113534
rect 6062 113298 6146 113534
rect 6382 113298 173094 113534
rect 173330 113298 173414 113534
rect 173650 113298 293826 113534
rect 294062 113298 294146 113534
rect 294382 113298 401826 113534
rect 402062 113298 402146 113534
rect 402382 113298 570350 113534
rect 570586 113298 570670 113534
rect 570906 113298 585342 113534
rect 585578 113298 585662 113534
rect 585898 113298 592650 113534
rect -8726 113266 592650 113298
rect -8726 82354 592650 82386
rect -8726 82118 -2934 82354
rect -2698 82118 -2614 82354
rect -2378 82118 13198 82354
rect 13434 82118 13518 82354
rect 13754 82118 167826 82354
rect 168062 82118 168146 82354
rect 168382 82118 291590 82354
rect 291826 82118 291910 82354
rect 292146 82118 419826 82354
rect 420062 82118 420146 82354
rect 420382 82118 563826 82354
rect 564062 82118 564146 82354
rect 564382 82118 582326 82354
rect 582562 82118 582646 82354
rect 582882 82118 586302 82354
rect 586538 82118 586622 82354
rect 586858 82118 592650 82354
rect -8726 82034 592650 82118
rect -8726 81798 -2934 82034
rect -2698 81798 -2614 82034
rect -2378 81798 13198 82034
rect 13434 81798 13518 82034
rect 13754 81798 167826 82034
rect 168062 81798 168146 82034
rect 168382 81798 291590 82034
rect 291826 81798 291910 82034
rect 292146 81798 419826 82034
rect 420062 81798 420146 82034
rect 420382 81798 563826 82034
rect 564062 81798 564146 82034
rect 564382 81798 582326 82034
rect 582562 81798 582646 82034
rect 582882 81798 586302 82034
rect 586538 81798 586622 82034
rect 586858 81798 592650 82034
rect -8726 81766 592650 81798
rect -8726 77854 592650 77886
rect -8726 77618 -1974 77854
rect -1738 77618 -1654 77854
rect -1418 77618 5826 77854
rect 6062 77618 6146 77854
rect 6382 77618 173094 77854
rect 173330 77618 173414 77854
rect 173650 77618 293826 77854
rect 294062 77618 294146 77854
rect 294382 77618 401826 77854
rect 402062 77618 402146 77854
rect 402382 77618 570350 77854
rect 570586 77618 570670 77854
rect 570906 77618 585342 77854
rect 585578 77618 585662 77854
rect 585898 77618 592650 77854
rect -8726 77534 592650 77618
rect -8726 77298 -1974 77534
rect -1738 77298 -1654 77534
rect -1418 77298 5826 77534
rect 6062 77298 6146 77534
rect 6382 77298 173094 77534
rect 173330 77298 173414 77534
rect 173650 77298 293826 77534
rect 294062 77298 294146 77534
rect 294382 77298 401826 77534
rect 402062 77298 402146 77534
rect 402382 77298 570350 77534
rect 570586 77298 570670 77534
rect 570906 77298 585342 77534
rect 585578 77298 585662 77534
rect 585898 77298 592650 77534
rect -8726 77266 592650 77298
rect -8726 46354 592650 46386
rect -8726 46118 -2934 46354
rect -2698 46118 -2614 46354
rect -2378 46118 13198 46354
rect 13434 46118 13518 46354
rect 13754 46118 167826 46354
rect 168062 46118 168146 46354
rect 168382 46118 291590 46354
rect 291826 46118 291910 46354
rect 292146 46118 419826 46354
rect 420062 46118 420146 46354
rect 420382 46118 563826 46354
rect 564062 46118 564146 46354
rect 564382 46118 582326 46354
rect 582562 46118 582646 46354
rect 582882 46118 586302 46354
rect 586538 46118 586622 46354
rect 586858 46118 592650 46354
rect -8726 46034 592650 46118
rect -8726 45798 -2934 46034
rect -2698 45798 -2614 46034
rect -2378 45798 13198 46034
rect 13434 45798 13518 46034
rect 13754 45798 167826 46034
rect 168062 45798 168146 46034
rect 168382 45798 291590 46034
rect 291826 45798 291910 46034
rect 292146 45798 419826 46034
rect 420062 45798 420146 46034
rect 420382 45798 563826 46034
rect 564062 45798 564146 46034
rect 564382 45798 582326 46034
rect 582562 45798 582646 46034
rect 582882 45798 586302 46034
rect 586538 45798 586622 46034
rect 586858 45798 592650 46034
rect -8726 45766 592650 45798
rect -8726 41854 592650 41886
rect -8726 41618 -1974 41854
rect -1738 41618 -1654 41854
rect -1418 41618 5826 41854
rect 6062 41618 6146 41854
rect 6382 41618 173094 41854
rect 173330 41618 173414 41854
rect 173650 41618 293826 41854
rect 294062 41618 294146 41854
rect 294382 41618 401826 41854
rect 402062 41618 402146 41854
rect 402382 41618 570350 41854
rect 570586 41618 570670 41854
rect 570906 41618 585342 41854
rect 585578 41618 585662 41854
rect 585898 41618 592650 41854
rect -8726 41534 592650 41618
rect -8726 41298 -1974 41534
rect -1738 41298 -1654 41534
rect -1418 41298 5826 41534
rect 6062 41298 6146 41534
rect 6382 41298 173094 41534
rect 173330 41298 173414 41534
rect 173650 41298 293826 41534
rect 294062 41298 294146 41534
rect 294382 41298 401826 41534
rect 402062 41298 402146 41534
rect 402382 41298 570350 41534
rect 570586 41298 570670 41534
rect 570906 41298 585342 41534
rect 585578 41298 585662 41534
rect 585898 41298 592650 41534
rect -8726 41266 592650 41298
rect -8726 10354 592650 10386
rect -8726 10118 -2934 10354
rect -2698 10118 -2614 10354
rect -2378 10118 23826 10354
rect 24062 10118 24146 10354
rect 24382 10118 59826 10354
rect 60062 10118 60146 10354
rect 60382 10118 95826 10354
rect 96062 10118 96146 10354
rect 96382 10118 131826 10354
rect 132062 10118 132146 10354
rect 132382 10118 167826 10354
rect 168062 10118 168146 10354
rect 168382 10118 203826 10354
rect 204062 10118 204146 10354
rect 204382 10118 239826 10354
rect 240062 10118 240146 10354
rect 240382 10118 275826 10354
rect 276062 10118 276146 10354
rect 276382 10118 311826 10354
rect 312062 10118 312146 10354
rect 312382 10118 347826 10354
rect 348062 10118 348146 10354
rect 348382 10118 383826 10354
rect 384062 10118 384146 10354
rect 384382 10118 419826 10354
rect 420062 10118 420146 10354
rect 420382 10118 455826 10354
rect 456062 10118 456146 10354
rect 456382 10118 491826 10354
rect 492062 10118 492146 10354
rect 492382 10118 527826 10354
rect 528062 10118 528146 10354
rect 528382 10118 563826 10354
rect 564062 10118 564146 10354
rect 564382 10118 582326 10354
rect 582562 10118 582646 10354
rect 582882 10118 586302 10354
rect 586538 10118 586622 10354
rect 586858 10118 592650 10354
rect -8726 10034 592650 10118
rect -8726 9798 -2934 10034
rect -2698 9798 -2614 10034
rect -2378 9798 23826 10034
rect 24062 9798 24146 10034
rect 24382 9798 59826 10034
rect 60062 9798 60146 10034
rect 60382 9798 95826 10034
rect 96062 9798 96146 10034
rect 96382 9798 131826 10034
rect 132062 9798 132146 10034
rect 132382 9798 167826 10034
rect 168062 9798 168146 10034
rect 168382 9798 203826 10034
rect 204062 9798 204146 10034
rect 204382 9798 239826 10034
rect 240062 9798 240146 10034
rect 240382 9798 275826 10034
rect 276062 9798 276146 10034
rect 276382 9798 311826 10034
rect 312062 9798 312146 10034
rect 312382 9798 347826 10034
rect 348062 9798 348146 10034
rect 348382 9798 383826 10034
rect 384062 9798 384146 10034
rect 384382 9798 419826 10034
rect 420062 9798 420146 10034
rect 420382 9798 455826 10034
rect 456062 9798 456146 10034
rect 456382 9798 491826 10034
rect 492062 9798 492146 10034
rect 492382 9798 527826 10034
rect 528062 9798 528146 10034
rect 528382 9798 563826 10034
rect 564062 9798 564146 10034
rect 564382 9798 582326 10034
rect 582562 9798 582646 10034
rect 582882 9798 586302 10034
rect 586538 9798 586622 10034
rect 586858 9798 592650 10034
rect -8726 9766 592650 9798
rect -8726 5854 592650 5886
rect -8726 5618 -1974 5854
rect -1738 5618 -1654 5854
rect -1418 5618 585342 5854
rect 585578 5618 585662 5854
rect 585898 5618 592650 5854
rect -8726 5534 592650 5618
rect -8726 5298 -1974 5534
rect -1738 5298 -1654 5534
rect -1418 5298 585342 5534
rect 585578 5298 585662 5534
rect 585898 5298 592650 5534
rect -8726 5266 592650 5298
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 582326 -1306
rect 582562 -1542 582646 -1306
rect 582882 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 582326 -1626
rect 582562 -1862 582646 -1626
rect 582882 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use Marmot  Marmot
timestamp 0
transform 1 0 4000 0 1 4000
box -960 -960 576960 696960
<< labels >>
flabel metal3 s 583520 285276 584960 285516 0 FreeSans 960 0 0 0 analog_io[0]
port 0 nsew signal bidirectional
flabel metal2 s 446098 703520 446210 704960 0 FreeSans 448 90 0 0 analog_io[10]
port 1 nsew signal bidirectional
flabel metal2 s 381146 703520 381258 704960 0 FreeSans 448 90 0 0 analog_io[11]
port 2 nsew signal bidirectional
flabel metal2 s 316286 703520 316398 704960 0 FreeSans 448 90 0 0 analog_io[12]
port 3 nsew signal bidirectional
flabel metal2 s 251426 703520 251538 704960 0 FreeSans 448 90 0 0 analog_io[13]
port 4 nsew signal bidirectional
flabel metal2 s 186474 703520 186586 704960 0 FreeSans 448 90 0 0 analog_io[14]
port 5 nsew signal bidirectional
flabel metal2 s 121614 703520 121726 704960 0 FreeSans 448 90 0 0 analog_io[15]
port 6 nsew signal bidirectional
flabel metal2 s 56754 703520 56866 704960 0 FreeSans 448 90 0 0 analog_io[16]
port 7 nsew signal bidirectional
flabel metal3 s -960 697220 480 697460 0 FreeSans 960 0 0 0 analog_io[17]
port 8 nsew signal bidirectional
flabel metal3 s -960 644996 480 645236 0 FreeSans 960 0 0 0 analog_io[18]
port 9 nsew signal bidirectional
flabel metal3 s -960 592908 480 593148 0 FreeSans 960 0 0 0 analog_io[19]
port 10 nsew signal bidirectional
flabel metal3 s 583520 338452 584960 338692 0 FreeSans 960 0 0 0 analog_io[1]
port 11 nsew signal bidirectional
flabel metal3 s -960 540684 480 540924 0 FreeSans 960 0 0 0 analog_io[20]
port 12 nsew signal bidirectional
flabel metal3 s -960 488596 480 488836 0 FreeSans 960 0 0 0 analog_io[21]
port 13 nsew signal bidirectional
flabel metal3 s -960 436508 480 436748 0 FreeSans 960 0 0 0 analog_io[22]
port 14 nsew signal bidirectional
flabel metal3 s -960 384284 480 384524 0 FreeSans 960 0 0 0 analog_io[23]
port 15 nsew signal bidirectional
flabel metal3 s -960 332196 480 332436 0 FreeSans 960 0 0 0 analog_io[24]
port 16 nsew signal bidirectional
flabel metal3 s -960 279972 480 280212 0 FreeSans 960 0 0 0 analog_io[25]
port 17 nsew signal bidirectional
flabel metal3 s -960 227884 480 228124 0 FreeSans 960 0 0 0 analog_io[26]
port 18 nsew signal bidirectional
flabel metal3 s -960 175796 480 176036 0 FreeSans 960 0 0 0 analog_io[27]
port 19 nsew signal bidirectional
flabel metal3 s -960 123572 480 123812 0 FreeSans 960 0 0 0 analog_io[28]
port 20 nsew signal bidirectional
flabel metal3 s 583520 391628 584960 391868 0 FreeSans 960 0 0 0 analog_io[2]
port 21 nsew signal bidirectional
flabel metal3 s 583520 444668 584960 444908 0 FreeSans 960 0 0 0 analog_io[3]
port 22 nsew signal bidirectional
flabel metal3 s 583520 497844 584960 498084 0 FreeSans 960 0 0 0 analog_io[4]
port 23 nsew signal bidirectional
flabel metal3 s 583520 551020 584960 551260 0 FreeSans 960 0 0 0 analog_io[5]
port 24 nsew signal bidirectional
flabel metal3 s 583520 604060 584960 604300 0 FreeSans 960 0 0 0 analog_io[6]
port 25 nsew signal bidirectional
flabel metal3 s 583520 657236 584960 657476 0 FreeSans 960 0 0 0 analog_io[7]
port 26 nsew signal bidirectional
flabel metal2 s 575818 703520 575930 704960 0 FreeSans 448 90 0 0 analog_io[8]
port 27 nsew signal bidirectional
flabel metal2 s 510958 703520 511070 704960 0 FreeSans 448 90 0 0 analog_io[9]
port 28 nsew signal bidirectional
flabel metal3 s 583520 6476 584960 6716 0 FreeSans 960 0 0 0 io_in[0]
port 29 nsew signal input
flabel metal3 s 583520 457996 584960 458236 0 FreeSans 960 0 0 0 io_in[10]
port 30 nsew signal input
flabel metal3 s 583520 511172 584960 511412 0 FreeSans 960 0 0 0 io_in[11]
port 31 nsew signal input
flabel metal3 s 583520 564212 584960 564452 0 FreeSans 960 0 0 0 io_in[12]
port 32 nsew signal input
flabel metal3 s 583520 617388 584960 617628 0 FreeSans 960 0 0 0 io_in[13]
port 33 nsew signal input
flabel metal3 s 583520 670564 584960 670804 0 FreeSans 960 0 0 0 io_in[14]
port 34 nsew signal input
flabel metal2 s 559626 703520 559738 704960 0 FreeSans 448 90 0 0 io_in[15]
port 35 nsew signal input
flabel metal2 s 494766 703520 494878 704960 0 FreeSans 448 90 0 0 io_in[16]
port 36 nsew signal input
flabel metal2 s 429814 703520 429926 704960 0 FreeSans 448 90 0 0 io_in[17]
port 37 nsew signal input
flabel metal2 s 364954 703520 365066 704960 0 FreeSans 448 90 0 0 io_in[18]
port 38 nsew signal input
flabel metal2 s 300094 703520 300206 704960 0 FreeSans 448 90 0 0 io_in[19]
port 39 nsew signal input
flabel metal3 s 583520 46188 584960 46428 0 FreeSans 960 0 0 0 io_in[1]
port 40 nsew signal input
flabel metal2 s 235142 703520 235254 704960 0 FreeSans 448 90 0 0 io_in[20]
port 41 nsew signal input
flabel metal2 s 170282 703520 170394 704960 0 FreeSans 448 90 0 0 io_in[21]
port 42 nsew signal input
flabel metal2 s 105422 703520 105534 704960 0 FreeSans 448 90 0 0 io_in[22]
port 43 nsew signal input
flabel metal2 s 40470 703520 40582 704960 0 FreeSans 448 90 0 0 io_in[23]
port 44 nsew signal input
flabel metal3 s -960 684164 480 684404 0 FreeSans 960 0 0 0 io_in[24]
port 45 nsew signal input
flabel metal3 s -960 631940 480 632180 0 FreeSans 960 0 0 0 io_in[25]
port 46 nsew signal input
flabel metal3 s -960 579852 480 580092 0 FreeSans 960 0 0 0 io_in[26]
port 47 nsew signal input
flabel metal3 s -960 527764 480 528004 0 FreeSans 960 0 0 0 io_in[27]
port 48 nsew signal input
flabel metal3 s -960 475540 480 475780 0 FreeSans 960 0 0 0 io_in[28]
port 49 nsew signal input
flabel metal3 s -960 423452 480 423692 0 FreeSans 960 0 0 0 io_in[29]
port 50 nsew signal input
flabel metal3 s 583520 86036 584960 86276 0 FreeSans 960 0 0 0 io_in[2]
port 51 nsew signal input
flabel metal3 s -960 371228 480 371468 0 FreeSans 960 0 0 0 io_in[30]
port 52 nsew signal input
flabel metal3 s -960 319140 480 319380 0 FreeSans 960 0 0 0 io_in[31]
port 53 nsew signal input
flabel metal3 s -960 267052 480 267292 0 FreeSans 960 0 0 0 io_in[32]
port 54 nsew signal input
flabel metal3 s -960 214828 480 215068 0 FreeSans 960 0 0 0 io_in[33]
port 55 nsew signal input
flabel metal3 s -960 162740 480 162980 0 FreeSans 960 0 0 0 io_in[34]
port 56 nsew signal input
flabel metal3 s -960 110516 480 110756 0 FreeSans 960 0 0 0 io_in[35]
port 57 nsew signal input
flabel metal3 s -960 71484 480 71724 0 FreeSans 960 0 0 0 io_in[36]
port 58 nsew signal input
flabel metal3 s -960 32316 480 32556 0 FreeSans 960 0 0 0 io_in[37]
port 59 nsew signal input
flabel metal3 s 583520 125884 584960 126124 0 FreeSans 960 0 0 0 io_in[3]
port 60 nsew signal input
flabel metal3 s 583520 165732 584960 165972 0 FreeSans 960 0 0 0 io_in[4]
port 61 nsew signal input
flabel metal3 s 583520 205580 584960 205820 0 FreeSans 960 0 0 0 io_in[5]
port 62 nsew signal input
flabel metal3 s 583520 245428 584960 245668 0 FreeSans 960 0 0 0 io_in[6]
port 63 nsew signal input
flabel metal3 s 583520 298604 584960 298844 0 FreeSans 960 0 0 0 io_in[7]
port 64 nsew signal input
flabel metal3 s 583520 351780 584960 352020 0 FreeSans 960 0 0 0 io_in[8]
port 65 nsew signal input
flabel metal3 s 583520 404820 584960 405060 0 FreeSans 960 0 0 0 io_in[9]
port 66 nsew signal input
flabel metal3 s 583520 32996 584960 33236 0 FreeSans 960 0 0 0 io_oeb[0]
port 67 nsew signal tristate
flabel metal3 s 583520 484516 584960 484756 0 FreeSans 960 0 0 0 io_oeb[10]
port 68 nsew signal tristate
flabel metal3 s 583520 537692 584960 537932 0 FreeSans 960 0 0 0 io_oeb[11]
port 69 nsew signal tristate
flabel metal3 s 583520 590868 584960 591108 0 FreeSans 960 0 0 0 io_oeb[12]
port 70 nsew signal tristate
flabel metal3 s 583520 643908 584960 644148 0 FreeSans 960 0 0 0 io_oeb[13]
port 71 nsew signal tristate
flabel metal3 s 583520 697084 584960 697324 0 FreeSans 960 0 0 0 io_oeb[14]
port 72 nsew signal tristate
flabel metal2 s 527150 703520 527262 704960 0 FreeSans 448 90 0 0 io_oeb[15]
port 73 nsew signal tristate
flabel metal2 s 462290 703520 462402 704960 0 FreeSans 448 90 0 0 io_oeb[16]
port 74 nsew signal tristate
flabel metal2 s 397430 703520 397542 704960 0 FreeSans 448 90 0 0 io_oeb[17]
port 75 nsew signal tristate
flabel metal2 s 332478 703520 332590 704960 0 FreeSans 448 90 0 0 io_oeb[18]
port 76 nsew signal tristate
flabel metal2 s 267618 703520 267730 704960 0 FreeSans 448 90 0 0 io_oeb[19]
port 77 nsew signal tristate
flabel metal3 s 583520 72844 584960 73084 0 FreeSans 960 0 0 0 io_oeb[1]
port 78 nsew signal tristate
flabel metal2 s 202758 703520 202870 704960 0 FreeSans 448 90 0 0 io_oeb[20]
port 79 nsew signal tristate
flabel metal2 s 137806 703520 137918 704960 0 FreeSans 448 90 0 0 io_oeb[21]
port 80 nsew signal tristate
flabel metal2 s 72946 703520 73058 704960 0 FreeSans 448 90 0 0 io_oeb[22]
port 81 nsew signal tristate
flabel metal2 s 8086 703520 8198 704960 0 FreeSans 448 90 0 0 io_oeb[23]
port 82 nsew signal tristate
flabel metal3 s -960 658052 480 658292 0 FreeSans 960 0 0 0 io_oeb[24]
port 83 nsew signal tristate
flabel metal3 s -960 605964 480 606204 0 FreeSans 960 0 0 0 io_oeb[25]
port 84 nsew signal tristate
flabel metal3 s -960 553740 480 553980 0 FreeSans 960 0 0 0 io_oeb[26]
port 85 nsew signal tristate
flabel metal3 s -960 501652 480 501892 0 FreeSans 960 0 0 0 io_oeb[27]
port 86 nsew signal tristate
flabel metal3 s -960 449428 480 449668 0 FreeSans 960 0 0 0 io_oeb[28]
port 87 nsew signal tristate
flabel metal3 s -960 397340 480 397580 0 FreeSans 960 0 0 0 io_oeb[29]
port 88 nsew signal tristate
flabel metal3 s 583520 112692 584960 112932 0 FreeSans 960 0 0 0 io_oeb[2]
port 89 nsew signal tristate
flabel metal3 s -960 345252 480 345492 0 FreeSans 960 0 0 0 io_oeb[30]
port 90 nsew signal tristate
flabel metal3 s -960 293028 480 293268 0 FreeSans 960 0 0 0 io_oeb[31]
port 91 nsew signal tristate
flabel metal3 s -960 240940 480 241180 0 FreeSans 960 0 0 0 io_oeb[32]
port 92 nsew signal tristate
flabel metal3 s -960 188716 480 188956 0 FreeSans 960 0 0 0 io_oeb[33]
port 93 nsew signal tristate
flabel metal3 s -960 136628 480 136868 0 FreeSans 960 0 0 0 io_oeb[34]
port 94 nsew signal tristate
flabel metal3 s -960 84540 480 84780 0 FreeSans 960 0 0 0 io_oeb[35]
port 95 nsew signal tristate
flabel metal3 s -960 45372 480 45612 0 FreeSans 960 0 0 0 io_oeb[36]
port 96 nsew signal tristate
flabel metal3 s -960 6340 480 6580 0 FreeSans 960 0 0 0 io_oeb[37]
port 97 nsew signal tristate
flabel metal3 s 583520 152540 584960 152780 0 FreeSans 960 0 0 0 io_oeb[3]
port 98 nsew signal tristate
flabel metal3 s 583520 192388 584960 192628 0 FreeSans 960 0 0 0 io_oeb[4]
port 99 nsew signal tristate
flabel metal3 s 583520 232236 584960 232476 0 FreeSans 960 0 0 0 io_oeb[5]
port 100 nsew signal tristate
flabel metal3 s 583520 272084 584960 272324 0 FreeSans 960 0 0 0 io_oeb[6]
port 101 nsew signal tristate
flabel metal3 s 583520 325124 584960 325364 0 FreeSans 960 0 0 0 io_oeb[7]
port 102 nsew signal tristate
flabel metal3 s 583520 378300 584960 378540 0 FreeSans 960 0 0 0 io_oeb[8]
port 103 nsew signal tristate
flabel metal3 s 583520 431476 584960 431716 0 FreeSans 960 0 0 0 io_oeb[9]
port 104 nsew signal tristate
flabel metal3 s 583520 19668 584960 19908 0 FreeSans 960 0 0 0 io_out[0]
port 105 nsew signal tristate
flabel metal3 s 583520 471324 584960 471564 0 FreeSans 960 0 0 0 io_out[10]
port 106 nsew signal tristate
flabel metal3 s 583520 524364 584960 524604 0 FreeSans 960 0 0 0 io_out[11]
port 107 nsew signal tristate
flabel metal3 s 583520 577540 584960 577780 0 FreeSans 960 0 0 0 io_out[12]
port 108 nsew signal tristate
flabel metal3 s 583520 630716 584960 630956 0 FreeSans 960 0 0 0 io_out[13]
port 109 nsew signal tristate
flabel metal3 s 583520 683756 584960 683996 0 FreeSans 960 0 0 0 io_out[14]
port 110 nsew signal tristate
flabel metal2 s 543434 703520 543546 704960 0 FreeSans 448 90 0 0 io_out[15]
port 111 nsew signal tristate
flabel metal2 s 478482 703520 478594 704960 0 FreeSans 448 90 0 0 io_out[16]
port 112 nsew signal tristate
flabel metal2 s 413622 703520 413734 704960 0 FreeSans 448 90 0 0 io_out[17]
port 113 nsew signal tristate
flabel metal2 s 348762 703520 348874 704960 0 FreeSans 448 90 0 0 io_out[18]
port 114 nsew signal tristate
flabel metal2 s 283810 703520 283922 704960 0 FreeSans 448 90 0 0 io_out[19]
port 115 nsew signal tristate
flabel metal3 s 583520 59516 584960 59756 0 FreeSans 960 0 0 0 io_out[1]
port 116 nsew signal tristate
flabel metal2 s 218950 703520 219062 704960 0 FreeSans 448 90 0 0 io_out[20]
port 117 nsew signal tristate
flabel metal2 s 154090 703520 154202 704960 0 FreeSans 448 90 0 0 io_out[21]
port 118 nsew signal tristate
flabel metal2 s 89138 703520 89250 704960 0 FreeSans 448 90 0 0 io_out[22]
port 119 nsew signal tristate
flabel metal2 s 24278 703520 24390 704960 0 FreeSans 448 90 0 0 io_out[23]
port 120 nsew signal tristate
flabel metal3 s -960 671108 480 671348 0 FreeSans 960 0 0 0 io_out[24]
port 121 nsew signal tristate
flabel metal3 s -960 619020 480 619260 0 FreeSans 960 0 0 0 io_out[25]
port 122 nsew signal tristate
flabel metal3 s -960 566796 480 567036 0 FreeSans 960 0 0 0 io_out[26]
port 123 nsew signal tristate
flabel metal3 s -960 514708 480 514948 0 FreeSans 960 0 0 0 io_out[27]
port 124 nsew signal tristate
flabel metal3 s -960 462484 480 462724 0 FreeSans 960 0 0 0 io_out[28]
port 125 nsew signal tristate
flabel metal3 s -960 410396 480 410636 0 FreeSans 960 0 0 0 io_out[29]
port 126 nsew signal tristate
flabel metal3 s 583520 99364 584960 99604 0 FreeSans 960 0 0 0 io_out[2]
port 127 nsew signal tristate
flabel metal3 s -960 358308 480 358548 0 FreeSans 960 0 0 0 io_out[30]
port 128 nsew signal tristate
flabel metal3 s -960 306084 480 306324 0 FreeSans 960 0 0 0 io_out[31]
port 129 nsew signal tristate
flabel metal3 s -960 253996 480 254236 0 FreeSans 960 0 0 0 io_out[32]
port 130 nsew signal tristate
flabel metal3 s -960 201772 480 202012 0 FreeSans 960 0 0 0 io_out[33]
port 131 nsew signal tristate
flabel metal3 s -960 149684 480 149924 0 FreeSans 960 0 0 0 io_out[34]
port 132 nsew signal tristate
flabel metal3 s -960 97460 480 97700 0 FreeSans 960 0 0 0 io_out[35]
port 133 nsew signal tristate
flabel metal3 s -960 58428 480 58668 0 FreeSans 960 0 0 0 io_out[36]
port 134 nsew signal tristate
flabel metal3 s -960 19260 480 19500 0 FreeSans 960 0 0 0 io_out[37]
port 135 nsew signal tristate
flabel metal3 s 583520 139212 584960 139452 0 FreeSans 960 0 0 0 io_out[3]
port 136 nsew signal tristate
flabel metal3 s 583520 179060 584960 179300 0 FreeSans 960 0 0 0 io_out[4]
port 137 nsew signal tristate
flabel metal3 s 583520 218908 584960 219148 0 FreeSans 960 0 0 0 io_out[5]
port 138 nsew signal tristate
flabel metal3 s 583520 258756 584960 258996 0 FreeSans 960 0 0 0 io_out[6]
port 139 nsew signal tristate
flabel metal3 s 583520 311932 584960 312172 0 FreeSans 960 0 0 0 io_out[7]
port 140 nsew signal tristate
flabel metal3 s 583520 364972 584960 365212 0 FreeSans 960 0 0 0 io_out[8]
port 141 nsew signal tristate
flabel metal3 s 583520 418148 584960 418388 0 FreeSans 960 0 0 0 io_out[9]
port 142 nsew signal tristate
flabel metal2 s 125846 -960 125958 480 0 FreeSans 448 90 0 0 la_data_in[0]
port 143 nsew signal input
flabel metal2 s 480506 -960 480618 480 0 FreeSans 448 90 0 0 la_data_in[100]
port 144 nsew signal input
flabel metal2 s 484002 -960 484114 480 0 FreeSans 448 90 0 0 la_data_in[101]
port 145 nsew signal input
flabel metal2 s 487590 -960 487702 480 0 FreeSans 448 90 0 0 la_data_in[102]
port 146 nsew signal input
flabel metal2 s 491086 -960 491198 480 0 FreeSans 448 90 0 0 la_data_in[103]
port 147 nsew signal input
flabel metal2 s 494674 -960 494786 480 0 FreeSans 448 90 0 0 la_data_in[104]
port 148 nsew signal input
flabel metal2 s 498170 -960 498282 480 0 FreeSans 448 90 0 0 la_data_in[105]
port 149 nsew signal input
flabel metal2 s 501758 -960 501870 480 0 FreeSans 448 90 0 0 la_data_in[106]
port 150 nsew signal input
flabel metal2 s 505346 -960 505458 480 0 FreeSans 448 90 0 0 la_data_in[107]
port 151 nsew signal input
flabel metal2 s 508842 -960 508954 480 0 FreeSans 448 90 0 0 la_data_in[108]
port 152 nsew signal input
flabel metal2 s 512430 -960 512542 480 0 FreeSans 448 90 0 0 la_data_in[109]
port 153 nsew signal input
flabel metal2 s 161266 -960 161378 480 0 FreeSans 448 90 0 0 la_data_in[10]
port 154 nsew signal input
flabel metal2 s 515926 -960 516038 480 0 FreeSans 448 90 0 0 la_data_in[110]
port 155 nsew signal input
flabel metal2 s 519514 -960 519626 480 0 FreeSans 448 90 0 0 la_data_in[111]
port 156 nsew signal input
flabel metal2 s 523010 -960 523122 480 0 FreeSans 448 90 0 0 la_data_in[112]
port 157 nsew signal input
flabel metal2 s 526598 -960 526710 480 0 FreeSans 448 90 0 0 la_data_in[113]
port 158 nsew signal input
flabel metal2 s 530094 -960 530206 480 0 FreeSans 448 90 0 0 la_data_in[114]
port 159 nsew signal input
flabel metal2 s 533682 -960 533794 480 0 FreeSans 448 90 0 0 la_data_in[115]
port 160 nsew signal input
flabel metal2 s 537178 -960 537290 480 0 FreeSans 448 90 0 0 la_data_in[116]
port 161 nsew signal input
flabel metal2 s 540766 -960 540878 480 0 FreeSans 448 90 0 0 la_data_in[117]
port 162 nsew signal input
flabel metal2 s 544354 -960 544466 480 0 FreeSans 448 90 0 0 la_data_in[118]
port 163 nsew signal input
flabel metal2 s 547850 -960 547962 480 0 FreeSans 448 90 0 0 la_data_in[119]
port 164 nsew signal input
flabel metal2 s 164854 -960 164966 480 0 FreeSans 448 90 0 0 la_data_in[11]
port 165 nsew signal input
flabel metal2 s 551438 -960 551550 480 0 FreeSans 448 90 0 0 la_data_in[120]
port 166 nsew signal input
flabel metal2 s 554934 -960 555046 480 0 FreeSans 448 90 0 0 la_data_in[121]
port 167 nsew signal input
flabel metal2 s 558522 -960 558634 480 0 FreeSans 448 90 0 0 la_data_in[122]
port 168 nsew signal input
flabel metal2 s 562018 -960 562130 480 0 FreeSans 448 90 0 0 la_data_in[123]
port 169 nsew signal input
flabel metal2 s 565606 -960 565718 480 0 FreeSans 448 90 0 0 la_data_in[124]
port 170 nsew signal input
flabel metal2 s 569102 -960 569214 480 0 FreeSans 448 90 0 0 la_data_in[125]
port 171 nsew signal input
flabel metal2 s 572690 -960 572802 480 0 FreeSans 448 90 0 0 la_data_in[126]
port 172 nsew signal input
flabel metal2 s 576278 -960 576390 480 0 FreeSans 448 90 0 0 la_data_in[127]
port 173 nsew signal input
flabel metal2 s 168350 -960 168462 480 0 FreeSans 448 90 0 0 la_data_in[12]
port 174 nsew signal input
flabel metal2 s 171938 -960 172050 480 0 FreeSans 448 90 0 0 la_data_in[13]
port 175 nsew signal input
flabel metal2 s 175434 -960 175546 480 0 FreeSans 448 90 0 0 la_data_in[14]
port 176 nsew signal input
flabel metal2 s 179022 -960 179134 480 0 FreeSans 448 90 0 0 la_data_in[15]
port 177 nsew signal input
flabel metal2 s 182518 -960 182630 480 0 FreeSans 448 90 0 0 la_data_in[16]
port 178 nsew signal input
flabel metal2 s 186106 -960 186218 480 0 FreeSans 448 90 0 0 la_data_in[17]
port 179 nsew signal input
flabel metal2 s 189694 -960 189806 480 0 FreeSans 448 90 0 0 la_data_in[18]
port 180 nsew signal input
flabel metal2 s 193190 -960 193302 480 0 FreeSans 448 90 0 0 la_data_in[19]
port 181 nsew signal input
flabel metal2 s 129342 -960 129454 480 0 FreeSans 448 90 0 0 la_data_in[1]
port 182 nsew signal input
flabel metal2 s 196778 -960 196890 480 0 FreeSans 448 90 0 0 la_data_in[20]
port 183 nsew signal input
flabel metal2 s 200274 -960 200386 480 0 FreeSans 448 90 0 0 la_data_in[21]
port 184 nsew signal input
flabel metal2 s 203862 -960 203974 480 0 FreeSans 448 90 0 0 la_data_in[22]
port 185 nsew signal input
flabel metal2 s 207358 -960 207470 480 0 FreeSans 448 90 0 0 la_data_in[23]
port 186 nsew signal input
flabel metal2 s 210946 -960 211058 480 0 FreeSans 448 90 0 0 la_data_in[24]
port 187 nsew signal input
flabel metal2 s 214442 -960 214554 480 0 FreeSans 448 90 0 0 la_data_in[25]
port 188 nsew signal input
flabel metal2 s 218030 -960 218142 480 0 FreeSans 448 90 0 0 la_data_in[26]
port 189 nsew signal input
flabel metal2 s 221526 -960 221638 480 0 FreeSans 448 90 0 0 la_data_in[27]
port 190 nsew signal input
flabel metal2 s 225114 -960 225226 480 0 FreeSans 448 90 0 0 la_data_in[28]
port 191 nsew signal input
flabel metal2 s 228702 -960 228814 480 0 FreeSans 448 90 0 0 la_data_in[29]
port 192 nsew signal input
flabel metal2 s 132930 -960 133042 480 0 FreeSans 448 90 0 0 la_data_in[2]
port 193 nsew signal input
flabel metal2 s 232198 -960 232310 480 0 FreeSans 448 90 0 0 la_data_in[30]
port 194 nsew signal input
flabel metal2 s 235786 -960 235898 480 0 FreeSans 448 90 0 0 la_data_in[31]
port 195 nsew signal input
flabel metal2 s 239282 -960 239394 480 0 FreeSans 448 90 0 0 la_data_in[32]
port 196 nsew signal input
flabel metal2 s 242870 -960 242982 480 0 FreeSans 448 90 0 0 la_data_in[33]
port 197 nsew signal input
flabel metal2 s 246366 -960 246478 480 0 FreeSans 448 90 0 0 la_data_in[34]
port 198 nsew signal input
flabel metal2 s 249954 -960 250066 480 0 FreeSans 448 90 0 0 la_data_in[35]
port 199 nsew signal input
flabel metal2 s 253450 -960 253562 480 0 FreeSans 448 90 0 0 la_data_in[36]
port 200 nsew signal input
flabel metal2 s 257038 -960 257150 480 0 FreeSans 448 90 0 0 la_data_in[37]
port 201 nsew signal input
flabel metal2 s 260626 -960 260738 480 0 FreeSans 448 90 0 0 la_data_in[38]
port 202 nsew signal input
flabel metal2 s 264122 -960 264234 480 0 FreeSans 448 90 0 0 la_data_in[39]
port 203 nsew signal input
flabel metal2 s 136426 -960 136538 480 0 FreeSans 448 90 0 0 la_data_in[3]
port 204 nsew signal input
flabel metal2 s 267710 -960 267822 480 0 FreeSans 448 90 0 0 la_data_in[40]
port 205 nsew signal input
flabel metal2 s 271206 -960 271318 480 0 FreeSans 448 90 0 0 la_data_in[41]
port 206 nsew signal input
flabel metal2 s 274794 -960 274906 480 0 FreeSans 448 90 0 0 la_data_in[42]
port 207 nsew signal input
flabel metal2 s 278290 -960 278402 480 0 FreeSans 448 90 0 0 la_data_in[43]
port 208 nsew signal input
flabel metal2 s 281878 -960 281990 480 0 FreeSans 448 90 0 0 la_data_in[44]
port 209 nsew signal input
flabel metal2 s 285374 -960 285486 480 0 FreeSans 448 90 0 0 la_data_in[45]
port 210 nsew signal input
flabel metal2 s 288962 -960 289074 480 0 FreeSans 448 90 0 0 la_data_in[46]
port 211 nsew signal input
flabel metal2 s 292550 -960 292662 480 0 FreeSans 448 90 0 0 la_data_in[47]
port 212 nsew signal input
flabel metal2 s 296046 -960 296158 480 0 FreeSans 448 90 0 0 la_data_in[48]
port 213 nsew signal input
flabel metal2 s 299634 -960 299746 480 0 FreeSans 448 90 0 0 la_data_in[49]
port 214 nsew signal input
flabel metal2 s 140014 -960 140126 480 0 FreeSans 448 90 0 0 la_data_in[4]
port 215 nsew signal input
flabel metal2 s 303130 -960 303242 480 0 FreeSans 448 90 0 0 la_data_in[50]
port 216 nsew signal input
flabel metal2 s 306718 -960 306830 480 0 FreeSans 448 90 0 0 la_data_in[51]
port 217 nsew signal input
flabel metal2 s 310214 -960 310326 480 0 FreeSans 448 90 0 0 la_data_in[52]
port 218 nsew signal input
flabel metal2 s 313802 -960 313914 480 0 FreeSans 448 90 0 0 la_data_in[53]
port 219 nsew signal input
flabel metal2 s 317298 -960 317410 480 0 FreeSans 448 90 0 0 la_data_in[54]
port 220 nsew signal input
flabel metal2 s 320886 -960 320998 480 0 FreeSans 448 90 0 0 la_data_in[55]
port 221 nsew signal input
flabel metal2 s 324382 -960 324494 480 0 FreeSans 448 90 0 0 la_data_in[56]
port 222 nsew signal input
flabel metal2 s 327970 -960 328082 480 0 FreeSans 448 90 0 0 la_data_in[57]
port 223 nsew signal input
flabel metal2 s 331558 -960 331670 480 0 FreeSans 448 90 0 0 la_data_in[58]
port 224 nsew signal input
flabel metal2 s 335054 -960 335166 480 0 FreeSans 448 90 0 0 la_data_in[59]
port 225 nsew signal input
flabel metal2 s 143510 -960 143622 480 0 FreeSans 448 90 0 0 la_data_in[5]
port 226 nsew signal input
flabel metal2 s 338642 -960 338754 480 0 FreeSans 448 90 0 0 la_data_in[60]
port 227 nsew signal input
flabel metal2 s 342138 -960 342250 480 0 FreeSans 448 90 0 0 la_data_in[61]
port 228 nsew signal input
flabel metal2 s 345726 -960 345838 480 0 FreeSans 448 90 0 0 la_data_in[62]
port 229 nsew signal input
flabel metal2 s 349222 -960 349334 480 0 FreeSans 448 90 0 0 la_data_in[63]
port 230 nsew signal input
flabel metal2 s 352810 -960 352922 480 0 FreeSans 448 90 0 0 la_data_in[64]
port 231 nsew signal input
flabel metal2 s 356306 -960 356418 480 0 FreeSans 448 90 0 0 la_data_in[65]
port 232 nsew signal input
flabel metal2 s 359894 -960 360006 480 0 FreeSans 448 90 0 0 la_data_in[66]
port 233 nsew signal input
flabel metal2 s 363482 -960 363594 480 0 FreeSans 448 90 0 0 la_data_in[67]
port 234 nsew signal input
flabel metal2 s 366978 -960 367090 480 0 FreeSans 448 90 0 0 la_data_in[68]
port 235 nsew signal input
flabel metal2 s 370566 -960 370678 480 0 FreeSans 448 90 0 0 la_data_in[69]
port 236 nsew signal input
flabel metal2 s 147098 -960 147210 480 0 FreeSans 448 90 0 0 la_data_in[6]
port 237 nsew signal input
flabel metal2 s 374062 -960 374174 480 0 FreeSans 448 90 0 0 la_data_in[70]
port 238 nsew signal input
flabel metal2 s 377650 -960 377762 480 0 FreeSans 448 90 0 0 la_data_in[71]
port 239 nsew signal input
flabel metal2 s 381146 -960 381258 480 0 FreeSans 448 90 0 0 la_data_in[72]
port 240 nsew signal input
flabel metal2 s 384734 -960 384846 480 0 FreeSans 448 90 0 0 la_data_in[73]
port 241 nsew signal input
flabel metal2 s 388230 -960 388342 480 0 FreeSans 448 90 0 0 la_data_in[74]
port 242 nsew signal input
flabel metal2 s 391818 -960 391930 480 0 FreeSans 448 90 0 0 la_data_in[75]
port 243 nsew signal input
flabel metal2 s 395314 -960 395426 480 0 FreeSans 448 90 0 0 la_data_in[76]
port 244 nsew signal input
flabel metal2 s 398902 -960 399014 480 0 FreeSans 448 90 0 0 la_data_in[77]
port 245 nsew signal input
flabel metal2 s 402490 -960 402602 480 0 FreeSans 448 90 0 0 la_data_in[78]
port 246 nsew signal input
flabel metal2 s 405986 -960 406098 480 0 FreeSans 448 90 0 0 la_data_in[79]
port 247 nsew signal input
flabel metal2 s 150594 -960 150706 480 0 FreeSans 448 90 0 0 la_data_in[7]
port 248 nsew signal input
flabel metal2 s 409574 -960 409686 480 0 FreeSans 448 90 0 0 la_data_in[80]
port 249 nsew signal input
flabel metal2 s 413070 -960 413182 480 0 FreeSans 448 90 0 0 la_data_in[81]
port 250 nsew signal input
flabel metal2 s 416658 -960 416770 480 0 FreeSans 448 90 0 0 la_data_in[82]
port 251 nsew signal input
flabel metal2 s 420154 -960 420266 480 0 FreeSans 448 90 0 0 la_data_in[83]
port 252 nsew signal input
flabel metal2 s 423742 -960 423854 480 0 FreeSans 448 90 0 0 la_data_in[84]
port 253 nsew signal input
flabel metal2 s 427238 -960 427350 480 0 FreeSans 448 90 0 0 la_data_in[85]
port 254 nsew signal input
flabel metal2 s 430826 -960 430938 480 0 FreeSans 448 90 0 0 la_data_in[86]
port 255 nsew signal input
flabel metal2 s 434414 -960 434526 480 0 FreeSans 448 90 0 0 la_data_in[87]
port 256 nsew signal input
flabel metal2 s 437910 -960 438022 480 0 FreeSans 448 90 0 0 la_data_in[88]
port 257 nsew signal input
flabel metal2 s 441498 -960 441610 480 0 FreeSans 448 90 0 0 la_data_in[89]
port 258 nsew signal input
flabel metal2 s 154182 -960 154294 480 0 FreeSans 448 90 0 0 la_data_in[8]
port 259 nsew signal input
flabel metal2 s 444994 -960 445106 480 0 FreeSans 448 90 0 0 la_data_in[90]
port 260 nsew signal input
flabel metal2 s 448582 -960 448694 480 0 FreeSans 448 90 0 0 la_data_in[91]
port 261 nsew signal input
flabel metal2 s 452078 -960 452190 480 0 FreeSans 448 90 0 0 la_data_in[92]
port 262 nsew signal input
flabel metal2 s 455666 -960 455778 480 0 FreeSans 448 90 0 0 la_data_in[93]
port 263 nsew signal input
flabel metal2 s 459162 -960 459274 480 0 FreeSans 448 90 0 0 la_data_in[94]
port 264 nsew signal input
flabel metal2 s 462750 -960 462862 480 0 FreeSans 448 90 0 0 la_data_in[95]
port 265 nsew signal input
flabel metal2 s 466246 -960 466358 480 0 FreeSans 448 90 0 0 la_data_in[96]
port 266 nsew signal input
flabel metal2 s 469834 -960 469946 480 0 FreeSans 448 90 0 0 la_data_in[97]
port 267 nsew signal input
flabel metal2 s 473422 -960 473534 480 0 FreeSans 448 90 0 0 la_data_in[98]
port 268 nsew signal input
flabel metal2 s 476918 -960 477030 480 0 FreeSans 448 90 0 0 la_data_in[99]
port 269 nsew signal input
flabel metal2 s 157770 -960 157882 480 0 FreeSans 448 90 0 0 la_data_in[9]
port 270 nsew signal input
flabel metal2 s 126950 -960 127062 480 0 FreeSans 448 90 0 0 la_data_out[0]
port 271 nsew signal tristate
flabel metal2 s 481702 -960 481814 480 0 FreeSans 448 90 0 0 la_data_out[100]
port 272 nsew signal tristate
flabel metal2 s 485198 -960 485310 480 0 FreeSans 448 90 0 0 la_data_out[101]
port 273 nsew signal tristate
flabel metal2 s 488786 -960 488898 480 0 FreeSans 448 90 0 0 la_data_out[102]
port 274 nsew signal tristate
flabel metal2 s 492282 -960 492394 480 0 FreeSans 448 90 0 0 la_data_out[103]
port 275 nsew signal tristate
flabel metal2 s 495870 -960 495982 480 0 FreeSans 448 90 0 0 la_data_out[104]
port 276 nsew signal tristate
flabel metal2 s 499366 -960 499478 480 0 FreeSans 448 90 0 0 la_data_out[105]
port 277 nsew signal tristate
flabel metal2 s 502954 -960 503066 480 0 FreeSans 448 90 0 0 la_data_out[106]
port 278 nsew signal tristate
flabel metal2 s 506450 -960 506562 480 0 FreeSans 448 90 0 0 la_data_out[107]
port 279 nsew signal tristate
flabel metal2 s 510038 -960 510150 480 0 FreeSans 448 90 0 0 la_data_out[108]
port 280 nsew signal tristate
flabel metal2 s 513534 -960 513646 480 0 FreeSans 448 90 0 0 la_data_out[109]
port 281 nsew signal tristate
flabel metal2 s 162462 -960 162574 480 0 FreeSans 448 90 0 0 la_data_out[10]
port 282 nsew signal tristate
flabel metal2 s 517122 -960 517234 480 0 FreeSans 448 90 0 0 la_data_out[110]
port 283 nsew signal tristate
flabel metal2 s 520710 -960 520822 480 0 FreeSans 448 90 0 0 la_data_out[111]
port 284 nsew signal tristate
flabel metal2 s 524206 -960 524318 480 0 FreeSans 448 90 0 0 la_data_out[112]
port 285 nsew signal tristate
flabel metal2 s 527794 -960 527906 480 0 FreeSans 448 90 0 0 la_data_out[113]
port 286 nsew signal tristate
flabel metal2 s 531290 -960 531402 480 0 FreeSans 448 90 0 0 la_data_out[114]
port 287 nsew signal tristate
flabel metal2 s 534878 -960 534990 480 0 FreeSans 448 90 0 0 la_data_out[115]
port 288 nsew signal tristate
flabel metal2 s 538374 -960 538486 480 0 FreeSans 448 90 0 0 la_data_out[116]
port 289 nsew signal tristate
flabel metal2 s 541962 -960 542074 480 0 FreeSans 448 90 0 0 la_data_out[117]
port 290 nsew signal tristate
flabel metal2 s 545458 -960 545570 480 0 FreeSans 448 90 0 0 la_data_out[118]
port 291 nsew signal tristate
flabel metal2 s 549046 -960 549158 480 0 FreeSans 448 90 0 0 la_data_out[119]
port 292 nsew signal tristate
flabel metal2 s 166050 -960 166162 480 0 FreeSans 448 90 0 0 la_data_out[11]
port 293 nsew signal tristate
flabel metal2 s 552634 -960 552746 480 0 FreeSans 448 90 0 0 la_data_out[120]
port 294 nsew signal tristate
flabel metal2 s 556130 -960 556242 480 0 FreeSans 448 90 0 0 la_data_out[121]
port 295 nsew signal tristate
flabel metal2 s 559718 -960 559830 480 0 FreeSans 448 90 0 0 la_data_out[122]
port 296 nsew signal tristate
flabel metal2 s 563214 -960 563326 480 0 FreeSans 448 90 0 0 la_data_out[123]
port 297 nsew signal tristate
flabel metal2 s 566802 -960 566914 480 0 FreeSans 448 90 0 0 la_data_out[124]
port 298 nsew signal tristate
flabel metal2 s 570298 -960 570410 480 0 FreeSans 448 90 0 0 la_data_out[125]
port 299 nsew signal tristate
flabel metal2 s 573886 -960 573998 480 0 FreeSans 448 90 0 0 la_data_out[126]
port 300 nsew signal tristate
flabel metal2 s 577382 -960 577494 480 0 FreeSans 448 90 0 0 la_data_out[127]
port 301 nsew signal tristate
flabel metal2 s 169546 -960 169658 480 0 FreeSans 448 90 0 0 la_data_out[12]
port 302 nsew signal tristate
flabel metal2 s 173134 -960 173246 480 0 FreeSans 448 90 0 0 la_data_out[13]
port 303 nsew signal tristate
flabel metal2 s 176630 -960 176742 480 0 FreeSans 448 90 0 0 la_data_out[14]
port 304 nsew signal tristate
flabel metal2 s 180218 -960 180330 480 0 FreeSans 448 90 0 0 la_data_out[15]
port 305 nsew signal tristate
flabel metal2 s 183714 -960 183826 480 0 FreeSans 448 90 0 0 la_data_out[16]
port 306 nsew signal tristate
flabel metal2 s 187302 -960 187414 480 0 FreeSans 448 90 0 0 la_data_out[17]
port 307 nsew signal tristate
flabel metal2 s 190798 -960 190910 480 0 FreeSans 448 90 0 0 la_data_out[18]
port 308 nsew signal tristate
flabel metal2 s 194386 -960 194498 480 0 FreeSans 448 90 0 0 la_data_out[19]
port 309 nsew signal tristate
flabel metal2 s 130538 -960 130650 480 0 FreeSans 448 90 0 0 la_data_out[1]
port 310 nsew signal tristate
flabel metal2 s 197882 -960 197994 480 0 FreeSans 448 90 0 0 la_data_out[20]
port 311 nsew signal tristate
flabel metal2 s 201470 -960 201582 480 0 FreeSans 448 90 0 0 la_data_out[21]
port 312 nsew signal tristate
flabel metal2 s 205058 -960 205170 480 0 FreeSans 448 90 0 0 la_data_out[22]
port 313 nsew signal tristate
flabel metal2 s 208554 -960 208666 480 0 FreeSans 448 90 0 0 la_data_out[23]
port 314 nsew signal tristate
flabel metal2 s 212142 -960 212254 480 0 FreeSans 448 90 0 0 la_data_out[24]
port 315 nsew signal tristate
flabel metal2 s 215638 -960 215750 480 0 FreeSans 448 90 0 0 la_data_out[25]
port 316 nsew signal tristate
flabel metal2 s 219226 -960 219338 480 0 FreeSans 448 90 0 0 la_data_out[26]
port 317 nsew signal tristate
flabel metal2 s 222722 -960 222834 480 0 FreeSans 448 90 0 0 la_data_out[27]
port 318 nsew signal tristate
flabel metal2 s 226310 -960 226422 480 0 FreeSans 448 90 0 0 la_data_out[28]
port 319 nsew signal tristate
flabel metal2 s 229806 -960 229918 480 0 FreeSans 448 90 0 0 la_data_out[29]
port 320 nsew signal tristate
flabel metal2 s 134126 -960 134238 480 0 FreeSans 448 90 0 0 la_data_out[2]
port 321 nsew signal tristate
flabel metal2 s 233394 -960 233506 480 0 FreeSans 448 90 0 0 la_data_out[30]
port 322 nsew signal tristate
flabel metal2 s 236982 -960 237094 480 0 FreeSans 448 90 0 0 la_data_out[31]
port 323 nsew signal tristate
flabel metal2 s 240478 -960 240590 480 0 FreeSans 448 90 0 0 la_data_out[32]
port 324 nsew signal tristate
flabel metal2 s 244066 -960 244178 480 0 FreeSans 448 90 0 0 la_data_out[33]
port 325 nsew signal tristate
flabel metal2 s 247562 -960 247674 480 0 FreeSans 448 90 0 0 la_data_out[34]
port 326 nsew signal tristate
flabel metal2 s 251150 -960 251262 480 0 FreeSans 448 90 0 0 la_data_out[35]
port 327 nsew signal tristate
flabel metal2 s 254646 -960 254758 480 0 FreeSans 448 90 0 0 la_data_out[36]
port 328 nsew signal tristate
flabel metal2 s 258234 -960 258346 480 0 FreeSans 448 90 0 0 la_data_out[37]
port 329 nsew signal tristate
flabel metal2 s 261730 -960 261842 480 0 FreeSans 448 90 0 0 la_data_out[38]
port 330 nsew signal tristate
flabel metal2 s 265318 -960 265430 480 0 FreeSans 448 90 0 0 la_data_out[39]
port 331 nsew signal tristate
flabel metal2 s 137622 -960 137734 480 0 FreeSans 448 90 0 0 la_data_out[3]
port 332 nsew signal tristate
flabel metal2 s 268814 -960 268926 480 0 FreeSans 448 90 0 0 la_data_out[40]
port 333 nsew signal tristate
flabel metal2 s 272402 -960 272514 480 0 FreeSans 448 90 0 0 la_data_out[41]
port 334 nsew signal tristate
flabel metal2 s 275990 -960 276102 480 0 FreeSans 448 90 0 0 la_data_out[42]
port 335 nsew signal tristate
flabel metal2 s 279486 -960 279598 480 0 FreeSans 448 90 0 0 la_data_out[43]
port 336 nsew signal tristate
flabel metal2 s 283074 -960 283186 480 0 FreeSans 448 90 0 0 la_data_out[44]
port 337 nsew signal tristate
flabel metal2 s 286570 -960 286682 480 0 FreeSans 448 90 0 0 la_data_out[45]
port 338 nsew signal tristate
flabel metal2 s 290158 -960 290270 480 0 FreeSans 448 90 0 0 la_data_out[46]
port 339 nsew signal tristate
flabel metal2 s 293654 -960 293766 480 0 FreeSans 448 90 0 0 la_data_out[47]
port 340 nsew signal tristate
flabel metal2 s 297242 -960 297354 480 0 FreeSans 448 90 0 0 la_data_out[48]
port 341 nsew signal tristate
flabel metal2 s 300738 -960 300850 480 0 FreeSans 448 90 0 0 la_data_out[49]
port 342 nsew signal tristate
flabel metal2 s 141210 -960 141322 480 0 FreeSans 448 90 0 0 la_data_out[4]
port 343 nsew signal tristate
flabel metal2 s 304326 -960 304438 480 0 FreeSans 448 90 0 0 la_data_out[50]
port 344 nsew signal tristate
flabel metal2 s 307914 -960 308026 480 0 FreeSans 448 90 0 0 la_data_out[51]
port 345 nsew signal tristate
flabel metal2 s 311410 -960 311522 480 0 FreeSans 448 90 0 0 la_data_out[52]
port 346 nsew signal tristate
flabel metal2 s 314998 -960 315110 480 0 FreeSans 448 90 0 0 la_data_out[53]
port 347 nsew signal tristate
flabel metal2 s 318494 -960 318606 480 0 FreeSans 448 90 0 0 la_data_out[54]
port 348 nsew signal tristate
flabel metal2 s 322082 -960 322194 480 0 FreeSans 448 90 0 0 la_data_out[55]
port 349 nsew signal tristate
flabel metal2 s 325578 -960 325690 480 0 FreeSans 448 90 0 0 la_data_out[56]
port 350 nsew signal tristate
flabel metal2 s 329166 -960 329278 480 0 FreeSans 448 90 0 0 la_data_out[57]
port 351 nsew signal tristate
flabel metal2 s 332662 -960 332774 480 0 FreeSans 448 90 0 0 la_data_out[58]
port 352 nsew signal tristate
flabel metal2 s 336250 -960 336362 480 0 FreeSans 448 90 0 0 la_data_out[59]
port 353 nsew signal tristate
flabel metal2 s 144706 -960 144818 480 0 FreeSans 448 90 0 0 la_data_out[5]
port 354 nsew signal tristate
flabel metal2 s 339838 -960 339950 480 0 FreeSans 448 90 0 0 la_data_out[60]
port 355 nsew signal tristate
flabel metal2 s 343334 -960 343446 480 0 FreeSans 448 90 0 0 la_data_out[61]
port 356 nsew signal tristate
flabel metal2 s 346922 -960 347034 480 0 FreeSans 448 90 0 0 la_data_out[62]
port 357 nsew signal tristate
flabel metal2 s 350418 -960 350530 480 0 FreeSans 448 90 0 0 la_data_out[63]
port 358 nsew signal tristate
flabel metal2 s 354006 -960 354118 480 0 FreeSans 448 90 0 0 la_data_out[64]
port 359 nsew signal tristate
flabel metal2 s 357502 -960 357614 480 0 FreeSans 448 90 0 0 la_data_out[65]
port 360 nsew signal tristate
flabel metal2 s 361090 -960 361202 480 0 FreeSans 448 90 0 0 la_data_out[66]
port 361 nsew signal tristate
flabel metal2 s 364586 -960 364698 480 0 FreeSans 448 90 0 0 la_data_out[67]
port 362 nsew signal tristate
flabel metal2 s 368174 -960 368286 480 0 FreeSans 448 90 0 0 la_data_out[68]
port 363 nsew signal tristate
flabel metal2 s 371670 -960 371782 480 0 FreeSans 448 90 0 0 la_data_out[69]
port 364 nsew signal tristate
flabel metal2 s 148294 -960 148406 480 0 FreeSans 448 90 0 0 la_data_out[6]
port 365 nsew signal tristate
flabel metal2 s 375258 -960 375370 480 0 FreeSans 448 90 0 0 la_data_out[70]
port 366 nsew signal tristate
flabel metal2 s 378846 -960 378958 480 0 FreeSans 448 90 0 0 la_data_out[71]
port 367 nsew signal tristate
flabel metal2 s 382342 -960 382454 480 0 FreeSans 448 90 0 0 la_data_out[72]
port 368 nsew signal tristate
flabel metal2 s 385930 -960 386042 480 0 FreeSans 448 90 0 0 la_data_out[73]
port 369 nsew signal tristate
flabel metal2 s 389426 -960 389538 480 0 FreeSans 448 90 0 0 la_data_out[74]
port 370 nsew signal tristate
flabel metal2 s 393014 -960 393126 480 0 FreeSans 448 90 0 0 la_data_out[75]
port 371 nsew signal tristate
flabel metal2 s 396510 -960 396622 480 0 FreeSans 448 90 0 0 la_data_out[76]
port 372 nsew signal tristate
flabel metal2 s 400098 -960 400210 480 0 FreeSans 448 90 0 0 la_data_out[77]
port 373 nsew signal tristate
flabel metal2 s 403594 -960 403706 480 0 FreeSans 448 90 0 0 la_data_out[78]
port 374 nsew signal tristate
flabel metal2 s 407182 -960 407294 480 0 FreeSans 448 90 0 0 la_data_out[79]
port 375 nsew signal tristate
flabel metal2 s 151790 -960 151902 480 0 FreeSans 448 90 0 0 la_data_out[7]
port 376 nsew signal tristate
flabel metal2 s 410770 -960 410882 480 0 FreeSans 448 90 0 0 la_data_out[80]
port 377 nsew signal tristate
flabel metal2 s 414266 -960 414378 480 0 FreeSans 448 90 0 0 la_data_out[81]
port 378 nsew signal tristate
flabel metal2 s 417854 -960 417966 480 0 FreeSans 448 90 0 0 la_data_out[82]
port 379 nsew signal tristate
flabel metal2 s 421350 -960 421462 480 0 FreeSans 448 90 0 0 la_data_out[83]
port 380 nsew signal tristate
flabel metal2 s 424938 -960 425050 480 0 FreeSans 448 90 0 0 la_data_out[84]
port 381 nsew signal tristate
flabel metal2 s 428434 -960 428546 480 0 FreeSans 448 90 0 0 la_data_out[85]
port 382 nsew signal tristate
flabel metal2 s 432022 -960 432134 480 0 FreeSans 448 90 0 0 la_data_out[86]
port 383 nsew signal tristate
flabel metal2 s 435518 -960 435630 480 0 FreeSans 448 90 0 0 la_data_out[87]
port 384 nsew signal tristate
flabel metal2 s 439106 -960 439218 480 0 FreeSans 448 90 0 0 la_data_out[88]
port 385 nsew signal tristate
flabel metal2 s 442602 -960 442714 480 0 FreeSans 448 90 0 0 la_data_out[89]
port 386 nsew signal tristate
flabel metal2 s 155378 -960 155490 480 0 FreeSans 448 90 0 0 la_data_out[8]
port 387 nsew signal tristate
flabel metal2 s 446190 -960 446302 480 0 FreeSans 448 90 0 0 la_data_out[90]
port 388 nsew signal tristate
flabel metal2 s 449778 -960 449890 480 0 FreeSans 448 90 0 0 la_data_out[91]
port 389 nsew signal tristate
flabel metal2 s 453274 -960 453386 480 0 FreeSans 448 90 0 0 la_data_out[92]
port 390 nsew signal tristate
flabel metal2 s 456862 -960 456974 480 0 FreeSans 448 90 0 0 la_data_out[93]
port 391 nsew signal tristate
flabel metal2 s 460358 -960 460470 480 0 FreeSans 448 90 0 0 la_data_out[94]
port 392 nsew signal tristate
flabel metal2 s 463946 -960 464058 480 0 FreeSans 448 90 0 0 la_data_out[95]
port 393 nsew signal tristate
flabel metal2 s 467442 -960 467554 480 0 FreeSans 448 90 0 0 la_data_out[96]
port 394 nsew signal tristate
flabel metal2 s 471030 -960 471142 480 0 FreeSans 448 90 0 0 la_data_out[97]
port 395 nsew signal tristate
flabel metal2 s 474526 -960 474638 480 0 FreeSans 448 90 0 0 la_data_out[98]
port 396 nsew signal tristate
flabel metal2 s 478114 -960 478226 480 0 FreeSans 448 90 0 0 la_data_out[99]
port 397 nsew signal tristate
flabel metal2 s 158874 -960 158986 480 0 FreeSans 448 90 0 0 la_data_out[9]
port 398 nsew signal tristate
flabel metal2 s 128146 -960 128258 480 0 FreeSans 448 90 0 0 la_oenb[0]
port 399 nsew signal input
flabel metal2 s 482806 -960 482918 480 0 FreeSans 448 90 0 0 la_oenb[100]
port 400 nsew signal input
flabel metal2 s 486394 -960 486506 480 0 FreeSans 448 90 0 0 la_oenb[101]
port 401 nsew signal input
flabel metal2 s 489890 -960 490002 480 0 FreeSans 448 90 0 0 la_oenb[102]
port 402 nsew signal input
flabel metal2 s 493478 -960 493590 480 0 FreeSans 448 90 0 0 la_oenb[103]
port 403 nsew signal input
flabel metal2 s 497066 -960 497178 480 0 FreeSans 448 90 0 0 la_oenb[104]
port 404 nsew signal input
flabel metal2 s 500562 -960 500674 480 0 FreeSans 448 90 0 0 la_oenb[105]
port 405 nsew signal input
flabel metal2 s 504150 -960 504262 480 0 FreeSans 448 90 0 0 la_oenb[106]
port 406 nsew signal input
flabel metal2 s 507646 -960 507758 480 0 FreeSans 448 90 0 0 la_oenb[107]
port 407 nsew signal input
flabel metal2 s 511234 -960 511346 480 0 FreeSans 448 90 0 0 la_oenb[108]
port 408 nsew signal input
flabel metal2 s 514730 -960 514842 480 0 FreeSans 448 90 0 0 la_oenb[109]
port 409 nsew signal input
flabel metal2 s 163658 -960 163770 480 0 FreeSans 448 90 0 0 la_oenb[10]
port 410 nsew signal input
flabel metal2 s 518318 -960 518430 480 0 FreeSans 448 90 0 0 la_oenb[110]
port 411 nsew signal input
flabel metal2 s 521814 -960 521926 480 0 FreeSans 448 90 0 0 la_oenb[111]
port 412 nsew signal input
flabel metal2 s 525402 -960 525514 480 0 FreeSans 448 90 0 0 la_oenb[112]
port 413 nsew signal input
flabel metal2 s 528990 -960 529102 480 0 FreeSans 448 90 0 0 la_oenb[113]
port 414 nsew signal input
flabel metal2 s 532486 -960 532598 480 0 FreeSans 448 90 0 0 la_oenb[114]
port 415 nsew signal input
flabel metal2 s 536074 -960 536186 480 0 FreeSans 448 90 0 0 la_oenb[115]
port 416 nsew signal input
flabel metal2 s 539570 -960 539682 480 0 FreeSans 448 90 0 0 la_oenb[116]
port 417 nsew signal input
flabel metal2 s 543158 -960 543270 480 0 FreeSans 448 90 0 0 la_oenb[117]
port 418 nsew signal input
flabel metal2 s 546654 -960 546766 480 0 FreeSans 448 90 0 0 la_oenb[118]
port 419 nsew signal input
flabel metal2 s 550242 -960 550354 480 0 FreeSans 448 90 0 0 la_oenb[119]
port 420 nsew signal input
flabel metal2 s 167154 -960 167266 480 0 FreeSans 448 90 0 0 la_oenb[11]
port 421 nsew signal input
flabel metal2 s 553738 -960 553850 480 0 FreeSans 448 90 0 0 la_oenb[120]
port 422 nsew signal input
flabel metal2 s 557326 -960 557438 480 0 FreeSans 448 90 0 0 la_oenb[121]
port 423 nsew signal input
flabel metal2 s 560822 -960 560934 480 0 FreeSans 448 90 0 0 la_oenb[122]
port 424 nsew signal input
flabel metal2 s 564410 -960 564522 480 0 FreeSans 448 90 0 0 la_oenb[123]
port 425 nsew signal input
flabel metal2 s 567998 -960 568110 480 0 FreeSans 448 90 0 0 la_oenb[124]
port 426 nsew signal input
flabel metal2 s 571494 -960 571606 480 0 FreeSans 448 90 0 0 la_oenb[125]
port 427 nsew signal input
flabel metal2 s 575082 -960 575194 480 0 FreeSans 448 90 0 0 la_oenb[126]
port 428 nsew signal input
flabel metal2 s 578578 -960 578690 480 0 FreeSans 448 90 0 0 la_oenb[127]
port 429 nsew signal input
flabel metal2 s 170742 -960 170854 480 0 FreeSans 448 90 0 0 la_oenb[12]
port 430 nsew signal input
flabel metal2 s 174238 -960 174350 480 0 FreeSans 448 90 0 0 la_oenb[13]
port 431 nsew signal input
flabel metal2 s 177826 -960 177938 480 0 FreeSans 448 90 0 0 la_oenb[14]
port 432 nsew signal input
flabel metal2 s 181414 -960 181526 480 0 FreeSans 448 90 0 0 la_oenb[15]
port 433 nsew signal input
flabel metal2 s 184910 -960 185022 480 0 FreeSans 448 90 0 0 la_oenb[16]
port 434 nsew signal input
flabel metal2 s 188498 -960 188610 480 0 FreeSans 448 90 0 0 la_oenb[17]
port 435 nsew signal input
flabel metal2 s 191994 -960 192106 480 0 FreeSans 448 90 0 0 la_oenb[18]
port 436 nsew signal input
flabel metal2 s 195582 -960 195694 480 0 FreeSans 448 90 0 0 la_oenb[19]
port 437 nsew signal input
flabel metal2 s 131734 -960 131846 480 0 FreeSans 448 90 0 0 la_oenb[1]
port 438 nsew signal input
flabel metal2 s 199078 -960 199190 480 0 FreeSans 448 90 0 0 la_oenb[20]
port 439 nsew signal input
flabel metal2 s 202666 -960 202778 480 0 FreeSans 448 90 0 0 la_oenb[21]
port 440 nsew signal input
flabel metal2 s 206162 -960 206274 480 0 FreeSans 448 90 0 0 la_oenb[22]
port 441 nsew signal input
flabel metal2 s 209750 -960 209862 480 0 FreeSans 448 90 0 0 la_oenb[23]
port 442 nsew signal input
flabel metal2 s 213338 -960 213450 480 0 FreeSans 448 90 0 0 la_oenb[24]
port 443 nsew signal input
flabel metal2 s 216834 -960 216946 480 0 FreeSans 448 90 0 0 la_oenb[25]
port 444 nsew signal input
flabel metal2 s 220422 -960 220534 480 0 FreeSans 448 90 0 0 la_oenb[26]
port 445 nsew signal input
flabel metal2 s 223918 -960 224030 480 0 FreeSans 448 90 0 0 la_oenb[27]
port 446 nsew signal input
flabel metal2 s 227506 -960 227618 480 0 FreeSans 448 90 0 0 la_oenb[28]
port 447 nsew signal input
flabel metal2 s 231002 -960 231114 480 0 FreeSans 448 90 0 0 la_oenb[29]
port 448 nsew signal input
flabel metal2 s 135230 -960 135342 480 0 FreeSans 448 90 0 0 la_oenb[2]
port 449 nsew signal input
flabel metal2 s 234590 -960 234702 480 0 FreeSans 448 90 0 0 la_oenb[30]
port 450 nsew signal input
flabel metal2 s 238086 -960 238198 480 0 FreeSans 448 90 0 0 la_oenb[31]
port 451 nsew signal input
flabel metal2 s 241674 -960 241786 480 0 FreeSans 448 90 0 0 la_oenb[32]
port 452 nsew signal input
flabel metal2 s 245170 -960 245282 480 0 FreeSans 448 90 0 0 la_oenb[33]
port 453 nsew signal input
flabel metal2 s 248758 -960 248870 480 0 FreeSans 448 90 0 0 la_oenb[34]
port 454 nsew signal input
flabel metal2 s 252346 -960 252458 480 0 FreeSans 448 90 0 0 la_oenb[35]
port 455 nsew signal input
flabel metal2 s 255842 -960 255954 480 0 FreeSans 448 90 0 0 la_oenb[36]
port 456 nsew signal input
flabel metal2 s 259430 -960 259542 480 0 FreeSans 448 90 0 0 la_oenb[37]
port 457 nsew signal input
flabel metal2 s 262926 -960 263038 480 0 FreeSans 448 90 0 0 la_oenb[38]
port 458 nsew signal input
flabel metal2 s 266514 -960 266626 480 0 FreeSans 448 90 0 0 la_oenb[39]
port 459 nsew signal input
flabel metal2 s 138818 -960 138930 480 0 FreeSans 448 90 0 0 la_oenb[3]
port 460 nsew signal input
flabel metal2 s 270010 -960 270122 480 0 FreeSans 448 90 0 0 la_oenb[40]
port 461 nsew signal input
flabel metal2 s 273598 -960 273710 480 0 FreeSans 448 90 0 0 la_oenb[41]
port 462 nsew signal input
flabel metal2 s 277094 -960 277206 480 0 FreeSans 448 90 0 0 la_oenb[42]
port 463 nsew signal input
flabel metal2 s 280682 -960 280794 480 0 FreeSans 448 90 0 0 la_oenb[43]
port 464 nsew signal input
flabel metal2 s 284270 -960 284382 480 0 FreeSans 448 90 0 0 la_oenb[44]
port 465 nsew signal input
flabel metal2 s 287766 -960 287878 480 0 FreeSans 448 90 0 0 la_oenb[45]
port 466 nsew signal input
flabel metal2 s 291354 -960 291466 480 0 FreeSans 448 90 0 0 la_oenb[46]
port 467 nsew signal input
flabel metal2 s 294850 -960 294962 480 0 FreeSans 448 90 0 0 la_oenb[47]
port 468 nsew signal input
flabel metal2 s 298438 -960 298550 480 0 FreeSans 448 90 0 0 la_oenb[48]
port 469 nsew signal input
flabel metal2 s 301934 -960 302046 480 0 FreeSans 448 90 0 0 la_oenb[49]
port 470 nsew signal input
flabel metal2 s 142406 -960 142518 480 0 FreeSans 448 90 0 0 la_oenb[4]
port 471 nsew signal input
flabel metal2 s 305522 -960 305634 480 0 FreeSans 448 90 0 0 la_oenb[50]
port 472 nsew signal input
flabel metal2 s 309018 -960 309130 480 0 FreeSans 448 90 0 0 la_oenb[51]
port 473 nsew signal input
flabel metal2 s 312606 -960 312718 480 0 FreeSans 448 90 0 0 la_oenb[52]
port 474 nsew signal input
flabel metal2 s 316194 -960 316306 480 0 FreeSans 448 90 0 0 la_oenb[53]
port 475 nsew signal input
flabel metal2 s 319690 -960 319802 480 0 FreeSans 448 90 0 0 la_oenb[54]
port 476 nsew signal input
flabel metal2 s 323278 -960 323390 480 0 FreeSans 448 90 0 0 la_oenb[55]
port 477 nsew signal input
flabel metal2 s 326774 -960 326886 480 0 FreeSans 448 90 0 0 la_oenb[56]
port 478 nsew signal input
flabel metal2 s 330362 -960 330474 480 0 FreeSans 448 90 0 0 la_oenb[57]
port 479 nsew signal input
flabel metal2 s 333858 -960 333970 480 0 FreeSans 448 90 0 0 la_oenb[58]
port 480 nsew signal input
flabel metal2 s 337446 -960 337558 480 0 FreeSans 448 90 0 0 la_oenb[59]
port 481 nsew signal input
flabel metal2 s 145902 -960 146014 480 0 FreeSans 448 90 0 0 la_oenb[5]
port 482 nsew signal input
flabel metal2 s 340942 -960 341054 480 0 FreeSans 448 90 0 0 la_oenb[60]
port 483 nsew signal input
flabel metal2 s 344530 -960 344642 480 0 FreeSans 448 90 0 0 la_oenb[61]
port 484 nsew signal input
flabel metal2 s 348026 -960 348138 480 0 FreeSans 448 90 0 0 la_oenb[62]
port 485 nsew signal input
flabel metal2 s 351614 -960 351726 480 0 FreeSans 448 90 0 0 la_oenb[63]
port 486 nsew signal input
flabel metal2 s 355202 -960 355314 480 0 FreeSans 448 90 0 0 la_oenb[64]
port 487 nsew signal input
flabel metal2 s 358698 -960 358810 480 0 FreeSans 448 90 0 0 la_oenb[65]
port 488 nsew signal input
flabel metal2 s 362286 -960 362398 480 0 FreeSans 448 90 0 0 la_oenb[66]
port 489 nsew signal input
flabel metal2 s 365782 -960 365894 480 0 FreeSans 448 90 0 0 la_oenb[67]
port 490 nsew signal input
flabel metal2 s 369370 -960 369482 480 0 FreeSans 448 90 0 0 la_oenb[68]
port 491 nsew signal input
flabel metal2 s 372866 -960 372978 480 0 FreeSans 448 90 0 0 la_oenb[69]
port 492 nsew signal input
flabel metal2 s 149490 -960 149602 480 0 FreeSans 448 90 0 0 la_oenb[6]
port 493 nsew signal input
flabel metal2 s 376454 -960 376566 480 0 FreeSans 448 90 0 0 la_oenb[70]
port 494 nsew signal input
flabel metal2 s 379950 -960 380062 480 0 FreeSans 448 90 0 0 la_oenb[71]
port 495 nsew signal input
flabel metal2 s 383538 -960 383650 480 0 FreeSans 448 90 0 0 la_oenb[72]
port 496 nsew signal input
flabel metal2 s 387126 -960 387238 480 0 FreeSans 448 90 0 0 la_oenb[73]
port 497 nsew signal input
flabel metal2 s 390622 -960 390734 480 0 FreeSans 448 90 0 0 la_oenb[74]
port 498 nsew signal input
flabel metal2 s 394210 -960 394322 480 0 FreeSans 448 90 0 0 la_oenb[75]
port 499 nsew signal input
flabel metal2 s 397706 -960 397818 480 0 FreeSans 448 90 0 0 la_oenb[76]
port 500 nsew signal input
flabel metal2 s 401294 -960 401406 480 0 FreeSans 448 90 0 0 la_oenb[77]
port 501 nsew signal input
flabel metal2 s 404790 -960 404902 480 0 FreeSans 448 90 0 0 la_oenb[78]
port 502 nsew signal input
flabel metal2 s 408378 -960 408490 480 0 FreeSans 448 90 0 0 la_oenb[79]
port 503 nsew signal input
flabel metal2 s 152986 -960 153098 480 0 FreeSans 448 90 0 0 la_oenb[7]
port 504 nsew signal input
flabel metal2 s 411874 -960 411986 480 0 FreeSans 448 90 0 0 la_oenb[80]
port 505 nsew signal input
flabel metal2 s 415462 -960 415574 480 0 FreeSans 448 90 0 0 la_oenb[81]
port 506 nsew signal input
flabel metal2 s 418958 -960 419070 480 0 FreeSans 448 90 0 0 la_oenb[82]
port 507 nsew signal input
flabel metal2 s 422546 -960 422658 480 0 FreeSans 448 90 0 0 la_oenb[83]
port 508 nsew signal input
flabel metal2 s 426134 -960 426246 480 0 FreeSans 448 90 0 0 la_oenb[84]
port 509 nsew signal input
flabel metal2 s 429630 -960 429742 480 0 FreeSans 448 90 0 0 la_oenb[85]
port 510 nsew signal input
flabel metal2 s 433218 -960 433330 480 0 FreeSans 448 90 0 0 la_oenb[86]
port 511 nsew signal input
flabel metal2 s 436714 -960 436826 480 0 FreeSans 448 90 0 0 la_oenb[87]
port 512 nsew signal input
flabel metal2 s 440302 -960 440414 480 0 FreeSans 448 90 0 0 la_oenb[88]
port 513 nsew signal input
flabel metal2 s 443798 -960 443910 480 0 FreeSans 448 90 0 0 la_oenb[89]
port 514 nsew signal input
flabel metal2 s 156574 -960 156686 480 0 FreeSans 448 90 0 0 la_oenb[8]
port 515 nsew signal input
flabel metal2 s 447386 -960 447498 480 0 FreeSans 448 90 0 0 la_oenb[90]
port 516 nsew signal input
flabel metal2 s 450882 -960 450994 480 0 FreeSans 448 90 0 0 la_oenb[91]
port 517 nsew signal input
flabel metal2 s 454470 -960 454582 480 0 FreeSans 448 90 0 0 la_oenb[92]
port 518 nsew signal input
flabel metal2 s 458058 -960 458170 480 0 FreeSans 448 90 0 0 la_oenb[93]
port 519 nsew signal input
flabel metal2 s 461554 -960 461666 480 0 FreeSans 448 90 0 0 la_oenb[94]
port 520 nsew signal input
flabel metal2 s 465142 -960 465254 480 0 FreeSans 448 90 0 0 la_oenb[95]
port 521 nsew signal input
flabel metal2 s 468638 -960 468750 480 0 FreeSans 448 90 0 0 la_oenb[96]
port 522 nsew signal input
flabel metal2 s 472226 -960 472338 480 0 FreeSans 448 90 0 0 la_oenb[97]
port 523 nsew signal input
flabel metal2 s 475722 -960 475834 480 0 FreeSans 448 90 0 0 la_oenb[98]
port 524 nsew signal input
flabel metal2 s 479310 -960 479422 480 0 FreeSans 448 90 0 0 la_oenb[99]
port 525 nsew signal input
flabel metal2 s 160070 -960 160182 480 0 FreeSans 448 90 0 0 la_oenb[9]
port 526 nsew signal input
flabel metal2 s 579774 -960 579886 480 0 FreeSans 448 90 0 0 user_clock2
port 527 nsew signal input
flabel metal2 s 580970 -960 581082 480 0 FreeSans 448 90 0 0 user_irq[0]
port 528 nsew signal tristate
flabel metal2 s 582166 -960 582278 480 0 FreeSans 448 90 0 0 user_irq[1]
port 529 nsew signal tristate
flabel metal2 s 583362 -960 583474 480 0 FreeSans 448 90 0 0 user_irq[2]
port 530 nsew signal tristate
flabel metal4 s -2006 -934 -1386 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 -934 585930 -314 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -2006 704250 585930 704870 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s 585310 -934 585930 704870 0 FreeSans 3840 90 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 5266 592650 5886 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 41266 592650 41886 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 77266 592650 77886 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 113266 592650 113886 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 149266 592650 149886 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 185266 592650 185886 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 221266 592650 221886 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 257266 592650 257886 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 293266 592650 293886 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 329266 592650 329886 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 365266 592650 365886 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 401266 592650 401886 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 437266 592650 437886 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 473266 592650 473886 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 509266 592650 509886 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 545266 592650 545886 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 581266 592650 581886 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 617266 592650 617886 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 653266 592650 653886 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal5 s -8726 689266 592650 689886 0 FreeSans 2560 0 0 0 vccd1
port 531 nsew power bidirectional
flabel metal4 s -3926 -2854 -3306 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 -2854 587850 -2234 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal5 s -3926 706170 587850 706790 0 FreeSans 2560 0 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s 587230 -2854 587850 706790 0 FreeSans 3840 90 0 0 vccd2
port 532 nsew power bidirectional
flabel metal4 s -5846 -4774 -5226 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 -4774 589770 -4154 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal5 s -5846 708090 589770 708710 0 FreeSans 2560 0 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s 589150 -4774 589770 708710 0 FreeSans 3840 90 0 0 vdda1
port 533 nsew power bidirectional
flabel metal4 s -7766 -6694 -7146 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 -6694 591690 -6074 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal5 s -7766 710010 591690 710630 0 FreeSans 2560 0 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s 591070 -6694 591690 710630 0 FreeSans 3840 90 0 0 vdda2
port 534 nsew power bidirectional
flabel metal4 s -6806 -5734 -6186 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 -5734 590730 -5114 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal5 s -6806 709050 590730 709670 0 FreeSans 2560 0 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s 590110 -5734 590730 709670 0 FreeSans 3840 90 0 0 vssa1
port 535 nsew ground bidirectional
flabel metal4 s -8726 -7654 -8106 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 -7654 592650 -7034 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal5 s -8726 710970 592650 711590 0 FreeSans 2560 0 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s 592030 -7654 592650 711590 0 FreeSans 3840 90 0 0 vssa2
port 536 nsew ground bidirectional
flabel metal4 s -2966 -1894 -2346 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 -1894 586890 -1274 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -2966 705210 586890 705830 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 586270 -1894 586890 705830 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s 582294 -7654 582914 711590 0 FreeSans 3840 90 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 9766 592650 10386 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 45766 592650 46386 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 81766 592650 82386 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 117766 592650 118386 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 153766 592650 154386 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 189766 592650 190386 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 225766 592650 226386 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 261766 592650 262386 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 297766 592650 298386 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 333766 592650 334386 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 369766 592650 370386 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 405766 592650 406386 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 441766 592650 442386 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 477766 592650 478386 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 513766 592650 514386 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 549766 592650 550386 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 585766 592650 586386 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 621766 592650 622386 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 657766 592650 658386 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal5 s -8726 693766 592650 694386 0 FreeSans 2560 0 0 0 vssd1
port 537 nsew ground bidirectional
flabel metal4 s -4886 -3814 -4266 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 -3814 588810 -3194 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal5 s -4886 707130 588810 707750 0 FreeSans 2560 0 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal4 s 588190 -3814 588810 707750 0 FreeSans 3840 90 0 0 vssd2
port 538 nsew ground bidirectional
flabel metal2 s 542 -960 654 480 0 FreeSans 448 90 0 0 wb_clk_i
port 539 nsew signal input
flabel metal2 s 1646 -960 1758 480 0 FreeSans 448 90 0 0 wb_rst_i
port 540 nsew signal input
flabel metal2 s 2842 -960 2954 480 0 FreeSans 448 90 0 0 wbs_ack_o
port 541 nsew signal tristate
flabel metal2 s 7626 -960 7738 480 0 FreeSans 448 90 0 0 wbs_adr_i[0]
port 542 nsew signal input
flabel metal2 s 47830 -960 47942 480 0 FreeSans 448 90 0 0 wbs_adr_i[10]
port 543 nsew signal input
flabel metal2 s 51326 -960 51438 480 0 FreeSans 448 90 0 0 wbs_adr_i[11]
port 544 nsew signal input
flabel metal2 s 54914 -960 55026 480 0 FreeSans 448 90 0 0 wbs_adr_i[12]
port 545 nsew signal input
flabel metal2 s 58410 -960 58522 480 0 FreeSans 448 90 0 0 wbs_adr_i[13]
port 546 nsew signal input
flabel metal2 s 61998 -960 62110 480 0 FreeSans 448 90 0 0 wbs_adr_i[14]
port 547 nsew signal input
flabel metal2 s 65494 -960 65606 480 0 FreeSans 448 90 0 0 wbs_adr_i[15]
port 548 nsew signal input
flabel metal2 s 69082 -960 69194 480 0 FreeSans 448 90 0 0 wbs_adr_i[16]
port 549 nsew signal input
flabel metal2 s 72578 -960 72690 480 0 FreeSans 448 90 0 0 wbs_adr_i[17]
port 550 nsew signal input
flabel metal2 s 76166 -960 76278 480 0 FreeSans 448 90 0 0 wbs_adr_i[18]
port 551 nsew signal input
flabel metal2 s 79662 -960 79774 480 0 FreeSans 448 90 0 0 wbs_adr_i[19]
port 552 nsew signal input
flabel metal2 s 12318 -960 12430 480 0 FreeSans 448 90 0 0 wbs_adr_i[1]
port 553 nsew signal input
flabel metal2 s 83250 -960 83362 480 0 FreeSans 448 90 0 0 wbs_adr_i[20]
port 554 nsew signal input
flabel metal2 s 86838 -960 86950 480 0 FreeSans 448 90 0 0 wbs_adr_i[21]
port 555 nsew signal input
flabel metal2 s 90334 -960 90446 480 0 FreeSans 448 90 0 0 wbs_adr_i[22]
port 556 nsew signal input
flabel metal2 s 93922 -960 94034 480 0 FreeSans 448 90 0 0 wbs_adr_i[23]
port 557 nsew signal input
flabel metal2 s 97418 -960 97530 480 0 FreeSans 448 90 0 0 wbs_adr_i[24]
port 558 nsew signal input
flabel metal2 s 101006 -960 101118 480 0 FreeSans 448 90 0 0 wbs_adr_i[25]
port 559 nsew signal input
flabel metal2 s 104502 -960 104614 480 0 FreeSans 448 90 0 0 wbs_adr_i[26]
port 560 nsew signal input
flabel metal2 s 108090 -960 108202 480 0 FreeSans 448 90 0 0 wbs_adr_i[27]
port 561 nsew signal input
flabel metal2 s 111586 -960 111698 480 0 FreeSans 448 90 0 0 wbs_adr_i[28]
port 562 nsew signal input
flabel metal2 s 115174 -960 115286 480 0 FreeSans 448 90 0 0 wbs_adr_i[29]
port 563 nsew signal input
flabel metal2 s 17010 -960 17122 480 0 FreeSans 448 90 0 0 wbs_adr_i[2]
port 564 nsew signal input
flabel metal2 s 118762 -960 118874 480 0 FreeSans 448 90 0 0 wbs_adr_i[30]
port 565 nsew signal input
flabel metal2 s 122258 -960 122370 480 0 FreeSans 448 90 0 0 wbs_adr_i[31]
port 566 nsew signal input
flabel metal2 s 21794 -960 21906 480 0 FreeSans 448 90 0 0 wbs_adr_i[3]
port 567 nsew signal input
flabel metal2 s 26486 -960 26598 480 0 FreeSans 448 90 0 0 wbs_adr_i[4]
port 568 nsew signal input
flabel metal2 s 30074 -960 30186 480 0 FreeSans 448 90 0 0 wbs_adr_i[5]
port 569 nsew signal input
flabel metal2 s 33570 -960 33682 480 0 FreeSans 448 90 0 0 wbs_adr_i[6]
port 570 nsew signal input
flabel metal2 s 37158 -960 37270 480 0 FreeSans 448 90 0 0 wbs_adr_i[7]
port 571 nsew signal input
flabel metal2 s 40654 -960 40766 480 0 FreeSans 448 90 0 0 wbs_adr_i[8]
port 572 nsew signal input
flabel metal2 s 44242 -960 44354 480 0 FreeSans 448 90 0 0 wbs_adr_i[9]
port 573 nsew signal input
flabel metal2 s 4038 -960 4150 480 0 FreeSans 448 90 0 0 wbs_cyc_i
port 574 nsew signal input
flabel metal2 s 8730 -960 8842 480 0 FreeSans 448 90 0 0 wbs_dat_i[0]
port 575 nsew signal input
flabel metal2 s 48934 -960 49046 480 0 FreeSans 448 90 0 0 wbs_dat_i[10]
port 576 nsew signal input
flabel metal2 s 52522 -960 52634 480 0 FreeSans 448 90 0 0 wbs_dat_i[11]
port 577 nsew signal input
flabel metal2 s 56018 -960 56130 480 0 FreeSans 448 90 0 0 wbs_dat_i[12]
port 578 nsew signal input
flabel metal2 s 59606 -960 59718 480 0 FreeSans 448 90 0 0 wbs_dat_i[13]
port 579 nsew signal input
flabel metal2 s 63194 -960 63306 480 0 FreeSans 448 90 0 0 wbs_dat_i[14]
port 580 nsew signal input
flabel metal2 s 66690 -960 66802 480 0 FreeSans 448 90 0 0 wbs_dat_i[15]
port 581 nsew signal input
flabel metal2 s 70278 -960 70390 480 0 FreeSans 448 90 0 0 wbs_dat_i[16]
port 582 nsew signal input
flabel metal2 s 73774 -960 73886 480 0 FreeSans 448 90 0 0 wbs_dat_i[17]
port 583 nsew signal input
flabel metal2 s 77362 -960 77474 480 0 FreeSans 448 90 0 0 wbs_dat_i[18]
port 584 nsew signal input
flabel metal2 s 80858 -960 80970 480 0 FreeSans 448 90 0 0 wbs_dat_i[19]
port 585 nsew signal input
flabel metal2 s 13514 -960 13626 480 0 FreeSans 448 90 0 0 wbs_dat_i[1]
port 586 nsew signal input
flabel metal2 s 84446 -960 84558 480 0 FreeSans 448 90 0 0 wbs_dat_i[20]
port 587 nsew signal input
flabel metal2 s 87942 -960 88054 480 0 FreeSans 448 90 0 0 wbs_dat_i[21]
port 588 nsew signal input
flabel metal2 s 91530 -960 91642 480 0 FreeSans 448 90 0 0 wbs_dat_i[22]
port 589 nsew signal input
flabel metal2 s 95118 -960 95230 480 0 FreeSans 448 90 0 0 wbs_dat_i[23]
port 590 nsew signal input
flabel metal2 s 98614 -960 98726 480 0 FreeSans 448 90 0 0 wbs_dat_i[24]
port 591 nsew signal input
flabel metal2 s 102202 -960 102314 480 0 FreeSans 448 90 0 0 wbs_dat_i[25]
port 592 nsew signal input
flabel metal2 s 105698 -960 105810 480 0 FreeSans 448 90 0 0 wbs_dat_i[26]
port 593 nsew signal input
flabel metal2 s 109286 -960 109398 480 0 FreeSans 448 90 0 0 wbs_dat_i[27]
port 594 nsew signal input
flabel metal2 s 112782 -960 112894 480 0 FreeSans 448 90 0 0 wbs_dat_i[28]
port 595 nsew signal input
flabel metal2 s 116370 -960 116482 480 0 FreeSans 448 90 0 0 wbs_dat_i[29]
port 596 nsew signal input
flabel metal2 s 18206 -960 18318 480 0 FreeSans 448 90 0 0 wbs_dat_i[2]
port 597 nsew signal input
flabel metal2 s 119866 -960 119978 480 0 FreeSans 448 90 0 0 wbs_dat_i[30]
port 598 nsew signal input
flabel metal2 s 123454 -960 123566 480 0 FreeSans 448 90 0 0 wbs_dat_i[31]
port 599 nsew signal input
flabel metal2 s 22990 -960 23102 480 0 FreeSans 448 90 0 0 wbs_dat_i[3]
port 600 nsew signal input
flabel metal2 s 27682 -960 27794 480 0 FreeSans 448 90 0 0 wbs_dat_i[4]
port 601 nsew signal input
flabel metal2 s 31270 -960 31382 480 0 FreeSans 448 90 0 0 wbs_dat_i[5]
port 602 nsew signal input
flabel metal2 s 34766 -960 34878 480 0 FreeSans 448 90 0 0 wbs_dat_i[6]
port 603 nsew signal input
flabel metal2 s 38354 -960 38466 480 0 FreeSans 448 90 0 0 wbs_dat_i[7]
port 604 nsew signal input
flabel metal2 s 41850 -960 41962 480 0 FreeSans 448 90 0 0 wbs_dat_i[8]
port 605 nsew signal input
flabel metal2 s 45438 -960 45550 480 0 FreeSans 448 90 0 0 wbs_dat_i[9]
port 606 nsew signal input
flabel metal2 s 9926 -960 10038 480 0 FreeSans 448 90 0 0 wbs_dat_o[0]
port 607 nsew signal tristate
flabel metal2 s 50130 -960 50242 480 0 FreeSans 448 90 0 0 wbs_dat_o[10]
port 608 nsew signal tristate
flabel metal2 s 53718 -960 53830 480 0 FreeSans 448 90 0 0 wbs_dat_o[11]
port 609 nsew signal tristate
flabel metal2 s 57214 -960 57326 480 0 FreeSans 448 90 0 0 wbs_dat_o[12]
port 610 nsew signal tristate
flabel metal2 s 60802 -960 60914 480 0 FreeSans 448 90 0 0 wbs_dat_o[13]
port 611 nsew signal tristate
flabel metal2 s 64298 -960 64410 480 0 FreeSans 448 90 0 0 wbs_dat_o[14]
port 612 nsew signal tristate
flabel metal2 s 67886 -960 67998 480 0 FreeSans 448 90 0 0 wbs_dat_o[15]
port 613 nsew signal tristate
flabel metal2 s 71474 -960 71586 480 0 FreeSans 448 90 0 0 wbs_dat_o[16]
port 614 nsew signal tristate
flabel metal2 s 74970 -960 75082 480 0 FreeSans 448 90 0 0 wbs_dat_o[17]
port 615 nsew signal tristate
flabel metal2 s 78558 -960 78670 480 0 FreeSans 448 90 0 0 wbs_dat_o[18]
port 616 nsew signal tristate
flabel metal2 s 82054 -960 82166 480 0 FreeSans 448 90 0 0 wbs_dat_o[19]
port 617 nsew signal tristate
flabel metal2 s 14710 -960 14822 480 0 FreeSans 448 90 0 0 wbs_dat_o[1]
port 618 nsew signal tristate
flabel metal2 s 85642 -960 85754 480 0 FreeSans 448 90 0 0 wbs_dat_o[20]
port 619 nsew signal tristate
flabel metal2 s 89138 -960 89250 480 0 FreeSans 448 90 0 0 wbs_dat_o[21]
port 620 nsew signal tristate
flabel metal2 s 92726 -960 92838 480 0 FreeSans 448 90 0 0 wbs_dat_o[22]
port 621 nsew signal tristate
flabel metal2 s 96222 -960 96334 480 0 FreeSans 448 90 0 0 wbs_dat_o[23]
port 622 nsew signal tristate
flabel metal2 s 99810 -960 99922 480 0 FreeSans 448 90 0 0 wbs_dat_o[24]
port 623 nsew signal tristate
flabel metal2 s 103306 -960 103418 480 0 FreeSans 448 90 0 0 wbs_dat_o[25]
port 624 nsew signal tristate
flabel metal2 s 106894 -960 107006 480 0 FreeSans 448 90 0 0 wbs_dat_o[26]
port 625 nsew signal tristate
flabel metal2 s 110482 -960 110594 480 0 FreeSans 448 90 0 0 wbs_dat_o[27]
port 626 nsew signal tristate
flabel metal2 s 113978 -960 114090 480 0 FreeSans 448 90 0 0 wbs_dat_o[28]
port 627 nsew signal tristate
flabel metal2 s 117566 -960 117678 480 0 FreeSans 448 90 0 0 wbs_dat_o[29]
port 628 nsew signal tristate
flabel metal2 s 19402 -960 19514 480 0 FreeSans 448 90 0 0 wbs_dat_o[2]
port 629 nsew signal tristate
flabel metal2 s 121062 -960 121174 480 0 FreeSans 448 90 0 0 wbs_dat_o[30]
port 630 nsew signal tristate
flabel metal2 s 124650 -960 124762 480 0 FreeSans 448 90 0 0 wbs_dat_o[31]
port 631 nsew signal tristate
flabel metal2 s 24186 -960 24298 480 0 FreeSans 448 90 0 0 wbs_dat_o[3]
port 632 nsew signal tristate
flabel metal2 s 28878 -960 28990 480 0 FreeSans 448 90 0 0 wbs_dat_o[4]
port 633 nsew signal tristate
flabel metal2 s 32374 -960 32486 480 0 FreeSans 448 90 0 0 wbs_dat_o[5]
port 634 nsew signal tristate
flabel metal2 s 35962 -960 36074 480 0 FreeSans 448 90 0 0 wbs_dat_o[6]
port 635 nsew signal tristate
flabel metal2 s 39550 -960 39662 480 0 FreeSans 448 90 0 0 wbs_dat_o[7]
port 636 nsew signal tristate
flabel metal2 s 43046 -960 43158 480 0 FreeSans 448 90 0 0 wbs_dat_o[8]
port 637 nsew signal tristate
flabel metal2 s 46634 -960 46746 480 0 FreeSans 448 90 0 0 wbs_dat_o[9]
port 638 nsew signal tristate
flabel metal2 s 11122 -960 11234 480 0 FreeSans 448 90 0 0 wbs_sel_i[0]
port 639 nsew signal input
flabel metal2 s 15906 -960 16018 480 0 FreeSans 448 90 0 0 wbs_sel_i[1]
port 640 nsew signal input
flabel metal2 s 20598 -960 20710 480 0 FreeSans 448 90 0 0 wbs_sel_i[2]
port 641 nsew signal input
flabel metal2 s 25290 -960 25402 480 0 FreeSans 448 90 0 0 wbs_sel_i[3]
port 642 nsew signal input
flabel metal2 s 5234 -960 5346 480 0 FreeSans 448 90 0 0 wbs_stb_i
port 643 nsew signal input
flabel metal2 s 6430 -960 6542 480 0 FreeSans 448 90 0 0 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
