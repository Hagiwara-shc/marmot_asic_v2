VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO Marmot
  CLASS BLOCK ;
  FOREIGN Marmot ;
  ORIGIN 0.000 0.000 ;
  SIZE 2880.000 BY 3480.000 ;
  PIN analog_io[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 1412.780 2884.800 1413.980 ;
    END
  END analog_io[0]
  PIN analog_io[10]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2195.530 3479.000 2196.090 3484.800 ;
    END
  END analog_io[10]
  PIN analog_io[11]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1877.210 3479.000 1877.770 3484.800 ;
    END
  END analog_io[11]
  PIN analog_io[12]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1558.890 3479.000 1559.450 3484.800 ;
    END
  END analog_io[12]
  PIN analog_io[13]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1240.570 3479.000 1241.130 3484.800 ;
    END
  END analog_io[13]
  PIN analog_io[14]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 922.250 3479.000 922.810 3484.800 ;
    END
  END analog_io[14]
  PIN analog_io[15]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 603.930 3479.000 604.490 3484.800 ;
    END
  END analog_io[15]
  PIN analog_io[16]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 285.610 3479.000 286.170 3484.800 ;
    END
  END analog_io[16]
  PIN analog_io[17]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3433.060 1.000 3434.260 ;
    END
  END analog_io[17]
  PIN analog_io[18]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3177.380 1.000 3178.580 ;
    END
  END analog_io[18]
  PIN analog_io[19]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2921.700 1.000 2922.900 ;
    END
  END analog_io[19]
  PIN analog_io[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 1673.900 2884.800 1675.100 ;
    END
  END analog_io[1]
  PIN analog_io[20]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2666.020 1.000 2667.220 ;
    END
  END analog_io[20]
  PIN analog_io[21]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2410.340 1.000 2411.540 ;
    END
  END analog_io[21]
  PIN analog_io[22]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2154.660 1.000 2155.860 ;
    END
  END analog_io[22]
  PIN analog_io[23]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1898.980 1.000 1900.180 ;
    END
  END analog_io[23]
  PIN analog_io[24]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1643.300 1.000 1644.500 ;
    END
  END analog_io[24]
  PIN analog_io[25]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1387.620 1.000 1388.820 ;
    END
  END analog_io[25]
  PIN analog_io[26]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1131.940 1.000 1133.140 ;
    END
  END analog_io[26]
  PIN analog_io[27]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 876.260 1.000 877.460 ;
    END
  END analog_io[27]
  PIN analog_io[28]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 620.580 1.000 621.780 ;
    END
  END analog_io[28]
  PIN analog_io[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 1935.020 2884.800 1936.220 ;
    END
  END analog_io[2]
  PIN analog_io[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 2196.140 2884.800 2197.340 ;
    END
  END analog_io[3]
  PIN analog_io[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 2457.260 2884.800 2458.460 ;
    END
  END analog_io[4]
  PIN analog_io[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 2718.380 2884.800 2719.580 ;
    END
  END analog_io[5]
  PIN analog_io[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 2979.500 2884.800 2980.700 ;
    END
  END analog_io[6]
  PIN analog_io[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 3240.620 2884.800 3241.820 ;
    END
  END analog_io[7]
  PIN analog_io[8]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2832.170 3479.000 2832.730 3484.800 ;
    END
  END analog_io[8]
  PIN analog_io[9]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2513.850 3479.000 2514.410 3484.800 ;
    END
  END analog_io[9]
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 41.900 2884.800 43.100 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 2261.420 2884.800 2262.620 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 2522.540 2884.800 2523.740 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 2783.660 2884.800 2784.860 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 3044.780 2884.800 3045.980 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 3305.900 2884.800 3307.100 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2752.590 3479.000 2753.150 3484.800 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2434.270 3479.000 2434.830 3484.800 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2115.950 3479.000 2116.510 3484.800 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1797.630 3479.000 1798.190 3484.800 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1479.310 3479.000 1479.870 3484.800 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 237.740 2884.800 238.940 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1160.990 3479.000 1161.550 3484.800 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 842.670 3479.000 843.230 3484.800 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 524.350 3479.000 524.910 3484.800 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 206.030 3479.000 206.590 3484.800 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3369.140 1.000 3370.340 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3113.460 1.000 3114.660 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2857.780 1.000 2858.980 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2602.100 1.000 2603.300 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2346.420 1.000 2347.620 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2090.740 1.000 2091.940 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 433.580 2884.800 434.780 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1835.060 1.000 1836.260 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1579.380 1.000 1580.580 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1323.700 1.000 1324.900 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1068.020 1.000 1069.220 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 812.340 1.000 813.540 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 556.660 1.000 557.860 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 364.900 1.000 366.100 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 173.140 1.000 174.340 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 629.420 2884.800 630.620 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 825.260 2884.800 826.460 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 1021.100 2884.800 1022.300 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 1216.940 2884.800 1218.140 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 1478.060 2884.800 1479.260 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 1739.180 2884.800 1740.380 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 2000.300 2884.800 2001.500 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 172.460 2884.800 173.660 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 2391.980 2884.800 2393.180 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 2653.100 2884.800 2654.300 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 2914.220 2884.800 2915.420 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 3175.340 2884.800 3176.540 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 3436.460 2884.800 3437.660 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2593.430 3479.000 2593.990 3484.800 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2275.110 3479.000 2275.670 3484.800 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1956.790 3479.000 1957.350 3484.800 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1638.470 3479.000 1639.030 3484.800 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1320.150 3479.000 1320.710 3484.800 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 368.300 2884.800 369.500 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1001.830 3479.000 1002.390 3484.800 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 683.510 3479.000 684.070 3484.800 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 365.190 3479.000 365.750 3484.800 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.870 3479.000 47.430 3484.800 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3241.300 1.000 3242.500 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2985.620 1.000 2986.820 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2729.940 1.000 2731.140 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2474.260 1.000 2475.460 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2218.580 1.000 2219.780 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1962.900 1.000 1964.100 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 564.140 2884.800 565.340 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1707.220 1.000 1708.420 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1451.540 1.000 1452.740 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1195.860 1.000 1197.060 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 940.180 1.000 941.380 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 684.500 1.000 685.700 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 428.820 1.000 430.020 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 237.060 1.000 238.260 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 45.300 1.000 46.500 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 759.980 2884.800 761.180 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 955.820 2884.800 957.020 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 1151.660 2884.800 1152.860 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 1347.500 2884.800 1348.700 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 1608.620 2884.800 1609.820 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 1869.740 2884.800 1870.940 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 2130.860 2884.800 2132.060 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 107.180 2884.800 108.380 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 2326.700 2884.800 2327.900 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 2587.820 2884.800 2589.020 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 2848.940 2884.800 2850.140 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 3110.060 2884.800 3111.260 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 3371.180 2884.800 3372.380 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2673.010 3479.000 2673.570 3484.800 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2354.690 3479.000 2355.250 3484.800 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2036.370 3479.000 2036.930 3484.800 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1718.050 3479.000 1718.610 3484.800 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1399.730 3479.000 1400.290 3484.800 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 303.020 2884.800 304.220 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1081.410 3479.000 1081.970 3484.800 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 763.090 3479.000 763.650 3484.800 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 444.770 3479.000 445.330 3484.800 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.450 3479.000 127.010 3484.800 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3305.220 1.000 3306.420 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 3049.540 1.000 3050.740 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2793.860 1.000 2795.060 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2538.180 1.000 2539.380 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2282.500 1.000 2283.700 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 2026.820 1.000 2028.020 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 498.860 2884.800 500.060 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1771.140 1.000 1772.340 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1515.460 1.000 1516.660 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1259.780 1.000 1260.980 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 1004.100 1.000 1005.300 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 748.420 1.000 749.620 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 492.740 1.000 493.940 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 300.980 1.000 302.180 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT -4.800 109.220 1.000 110.420 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 694.700 2884.800 695.900 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 890.540 2884.800 891.740 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 1086.380 2884.800 1087.580 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 1282.220 2884.800 1283.420 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 1543.340 2884.800 1544.540 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 1804.460 2884.800 1805.660 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 2879.000 2065.580 2884.800 2066.780 ;
    END
  END io_out[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 664.190 -4.800 664.750 1.000 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2320.190 -4.800 2320.750 1.000 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2336.750 -4.800 2337.310 1.000 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2353.310 -4.800 2353.870 1.000 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2369.870 -4.800 2370.430 1.000 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2386.430 -4.800 2386.990 1.000 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2402.990 -4.800 2403.550 1.000 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2419.550 -4.800 2420.110 1.000 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2436.110 -4.800 2436.670 1.000 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2452.670 -4.800 2453.230 1.000 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2469.230 -4.800 2469.790 1.000 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 829.790 -4.800 830.350 1.000 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2485.790 -4.800 2486.350 1.000 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2502.350 -4.800 2502.910 1.000 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2518.910 -4.800 2519.470 1.000 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2535.470 -4.800 2536.030 1.000 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2552.030 -4.800 2552.590 1.000 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2568.590 -4.800 2569.150 1.000 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2585.150 -4.800 2585.710 1.000 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2601.710 -4.800 2602.270 1.000 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2618.270 -4.800 2618.830 1.000 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2634.830 -4.800 2635.390 1.000 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 846.350 -4.800 846.910 1.000 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2651.390 -4.800 2651.950 1.000 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2667.950 -4.800 2668.510 1.000 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2684.510 -4.800 2685.070 1.000 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2701.070 -4.800 2701.630 1.000 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2717.630 -4.800 2718.190 1.000 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2734.190 -4.800 2734.750 1.000 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2750.750 -4.800 2751.310 1.000 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2767.310 -4.800 2767.870 1.000 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 862.910 -4.800 863.470 1.000 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 879.470 -4.800 880.030 1.000 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 896.030 -4.800 896.590 1.000 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 912.590 -4.800 913.150 1.000 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 929.150 -4.800 929.710 1.000 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 945.710 -4.800 946.270 1.000 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 962.270 -4.800 962.830 1.000 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 978.830 -4.800 979.390 1.000 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 680.750 -4.800 681.310 1.000 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 995.390 -4.800 995.950 1.000 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1011.950 -4.800 1012.510 1.000 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1028.510 -4.800 1029.070 1.000 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1045.070 -4.800 1045.630 1.000 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1061.630 -4.800 1062.190 1.000 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1078.190 -4.800 1078.750 1.000 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1094.750 -4.800 1095.310 1.000 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1111.310 -4.800 1111.870 1.000 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1127.870 -4.800 1128.430 1.000 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1144.430 -4.800 1144.990 1.000 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 697.310 -4.800 697.870 1.000 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1160.990 -4.800 1161.550 1.000 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1177.550 -4.800 1178.110 1.000 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1194.110 -4.800 1194.670 1.000 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1210.670 -4.800 1211.230 1.000 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1227.230 -4.800 1227.790 1.000 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1243.790 -4.800 1244.350 1.000 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1260.350 -4.800 1260.910 1.000 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1276.910 -4.800 1277.470 1.000 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1293.470 -4.800 1294.030 1.000 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1310.030 -4.800 1310.590 1.000 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 713.870 -4.800 714.430 1.000 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1326.590 -4.800 1327.150 1.000 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1343.150 -4.800 1343.710 1.000 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1359.710 -4.800 1360.270 1.000 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1376.270 -4.800 1376.830 1.000 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1392.830 -4.800 1393.390 1.000 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1409.390 -4.800 1409.950 1.000 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1425.950 -4.800 1426.510 1.000 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1442.510 -4.800 1443.070 1.000 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1459.070 -4.800 1459.630 1.000 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1475.630 -4.800 1476.190 1.000 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 730.430 -4.800 730.990 1.000 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1492.190 -4.800 1492.750 1.000 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1508.750 -4.800 1509.310 1.000 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1525.310 -4.800 1525.870 1.000 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1541.870 -4.800 1542.430 1.000 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1558.430 -4.800 1558.990 1.000 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1574.990 -4.800 1575.550 1.000 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1591.550 -4.800 1592.110 1.000 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1608.110 -4.800 1608.670 1.000 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1624.670 -4.800 1625.230 1.000 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1641.230 -4.800 1641.790 1.000 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 746.990 -4.800 747.550 1.000 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1657.790 -4.800 1658.350 1.000 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1674.350 -4.800 1674.910 1.000 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1690.910 -4.800 1691.470 1.000 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1707.470 -4.800 1708.030 1.000 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1724.030 -4.800 1724.590 1.000 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1740.590 -4.800 1741.150 1.000 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1757.150 -4.800 1757.710 1.000 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1773.710 -4.800 1774.270 1.000 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1790.270 -4.800 1790.830 1.000 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1806.830 -4.800 1807.390 1.000 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 763.550 -4.800 764.110 1.000 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1823.390 -4.800 1823.950 1.000 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1839.950 -4.800 1840.510 1.000 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1856.510 -4.800 1857.070 1.000 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1873.070 -4.800 1873.630 1.000 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1889.630 -4.800 1890.190 1.000 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1906.190 -4.800 1906.750 1.000 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1922.750 -4.800 1923.310 1.000 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1939.310 -4.800 1939.870 1.000 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1955.870 -4.800 1956.430 1.000 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1972.430 -4.800 1972.990 1.000 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 780.110 -4.800 780.670 1.000 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1988.990 -4.800 1989.550 1.000 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2005.550 -4.800 2006.110 1.000 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2022.110 -4.800 2022.670 1.000 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2038.670 -4.800 2039.230 1.000 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2055.230 -4.800 2055.790 1.000 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2071.790 -4.800 2072.350 1.000 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2088.350 -4.800 2088.910 1.000 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2104.910 -4.800 2105.470 1.000 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2121.470 -4.800 2122.030 1.000 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2138.030 -4.800 2138.590 1.000 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 796.670 -4.800 797.230 1.000 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2154.590 -4.800 2155.150 1.000 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2171.150 -4.800 2171.710 1.000 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2187.710 -4.800 2188.270 1.000 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2204.270 -4.800 2204.830 1.000 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2220.830 -4.800 2221.390 1.000 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2237.390 -4.800 2237.950 1.000 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2253.950 -4.800 2254.510 1.000 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2270.510 -4.800 2271.070 1.000 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2287.070 -4.800 2287.630 1.000 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2303.630 -4.800 2304.190 1.000 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 813.230 -4.800 813.790 1.000 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 669.710 -4.800 670.270 1.000 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2325.710 -4.800 2326.270 1.000 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2342.270 -4.800 2342.830 1.000 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2358.830 -4.800 2359.390 1.000 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2375.390 -4.800 2375.950 1.000 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2391.950 -4.800 2392.510 1.000 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2408.510 -4.800 2409.070 1.000 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2425.070 -4.800 2425.630 1.000 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2441.630 -4.800 2442.190 1.000 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2458.190 -4.800 2458.750 1.000 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2474.750 -4.800 2475.310 1.000 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 835.310 -4.800 835.870 1.000 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2491.310 -4.800 2491.870 1.000 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2507.870 -4.800 2508.430 1.000 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2524.430 -4.800 2524.990 1.000 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2540.990 -4.800 2541.550 1.000 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2557.550 -4.800 2558.110 1.000 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2574.110 -4.800 2574.670 1.000 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2590.670 -4.800 2591.230 1.000 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2607.230 -4.800 2607.790 1.000 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2623.790 -4.800 2624.350 1.000 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2640.350 -4.800 2640.910 1.000 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 851.870 -4.800 852.430 1.000 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2656.910 -4.800 2657.470 1.000 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2673.470 -4.800 2674.030 1.000 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2690.030 -4.800 2690.590 1.000 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2706.590 -4.800 2707.150 1.000 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2723.150 -4.800 2723.710 1.000 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2739.710 -4.800 2740.270 1.000 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2756.270 -4.800 2756.830 1.000 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2772.830 -4.800 2773.390 1.000 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 868.430 -4.800 868.990 1.000 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 884.990 -4.800 885.550 1.000 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 901.550 -4.800 902.110 1.000 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 918.110 -4.800 918.670 1.000 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 934.670 -4.800 935.230 1.000 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 951.230 -4.800 951.790 1.000 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 967.790 -4.800 968.350 1.000 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 984.350 -4.800 984.910 1.000 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 686.270 -4.800 686.830 1.000 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1000.910 -4.800 1001.470 1.000 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1017.470 -4.800 1018.030 1.000 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1034.030 -4.800 1034.590 1.000 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1050.590 -4.800 1051.150 1.000 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1067.150 -4.800 1067.710 1.000 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1083.710 -4.800 1084.270 1.000 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1100.270 -4.800 1100.830 1.000 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1116.830 -4.800 1117.390 1.000 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1133.390 -4.800 1133.950 1.000 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1149.950 -4.800 1150.510 1.000 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 702.830 -4.800 703.390 1.000 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1166.510 -4.800 1167.070 1.000 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1183.070 -4.800 1183.630 1.000 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1199.630 -4.800 1200.190 1.000 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1216.190 -4.800 1216.750 1.000 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1232.750 -4.800 1233.310 1.000 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1249.310 -4.800 1249.870 1.000 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1265.870 -4.800 1266.430 1.000 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1282.430 -4.800 1282.990 1.000 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1298.990 -4.800 1299.550 1.000 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1315.550 -4.800 1316.110 1.000 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 719.390 -4.800 719.950 1.000 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1332.110 -4.800 1332.670 1.000 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1348.670 -4.800 1349.230 1.000 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1365.230 -4.800 1365.790 1.000 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1381.790 -4.800 1382.350 1.000 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1398.350 -4.800 1398.910 1.000 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1414.910 -4.800 1415.470 1.000 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1431.470 -4.800 1432.030 1.000 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1448.030 -4.800 1448.590 1.000 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1464.590 -4.800 1465.150 1.000 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1481.150 -4.800 1481.710 1.000 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 735.950 -4.800 736.510 1.000 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1497.710 -4.800 1498.270 1.000 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1514.270 -4.800 1514.830 1.000 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1530.830 -4.800 1531.390 1.000 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1547.390 -4.800 1547.950 1.000 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1563.950 -4.800 1564.510 1.000 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1580.510 -4.800 1581.070 1.000 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1597.070 -4.800 1597.630 1.000 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1613.630 -4.800 1614.190 1.000 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1630.190 -4.800 1630.750 1.000 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1646.750 -4.800 1647.310 1.000 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 752.510 -4.800 753.070 1.000 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1663.310 -4.800 1663.870 1.000 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1679.870 -4.800 1680.430 1.000 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1696.430 -4.800 1696.990 1.000 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1712.990 -4.800 1713.550 1.000 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1729.550 -4.800 1730.110 1.000 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1746.110 -4.800 1746.670 1.000 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1762.670 -4.800 1763.230 1.000 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1779.230 -4.800 1779.790 1.000 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1795.790 -4.800 1796.350 1.000 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1812.350 -4.800 1812.910 1.000 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 769.070 -4.800 769.630 1.000 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1828.910 -4.800 1829.470 1.000 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1845.470 -4.800 1846.030 1.000 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1862.030 -4.800 1862.590 1.000 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1878.590 -4.800 1879.150 1.000 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1895.150 -4.800 1895.710 1.000 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1911.710 -4.800 1912.270 1.000 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1928.270 -4.800 1928.830 1.000 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1944.830 -4.800 1945.390 1.000 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1961.390 -4.800 1961.950 1.000 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1977.950 -4.800 1978.510 1.000 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 785.630 -4.800 786.190 1.000 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1994.510 -4.800 1995.070 1.000 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2011.070 -4.800 2011.630 1.000 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2027.630 -4.800 2028.190 1.000 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2044.190 -4.800 2044.750 1.000 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2060.750 -4.800 2061.310 1.000 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2077.310 -4.800 2077.870 1.000 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2093.870 -4.800 2094.430 1.000 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2110.430 -4.800 2110.990 1.000 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2126.990 -4.800 2127.550 1.000 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2143.550 -4.800 2144.110 1.000 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 802.190 -4.800 802.750 1.000 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2160.110 -4.800 2160.670 1.000 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2176.670 -4.800 2177.230 1.000 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2193.230 -4.800 2193.790 1.000 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2209.790 -4.800 2210.350 1.000 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2226.350 -4.800 2226.910 1.000 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2242.910 -4.800 2243.470 1.000 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2259.470 -4.800 2260.030 1.000 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2276.030 -4.800 2276.590 1.000 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2292.590 -4.800 2293.150 1.000 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2309.150 -4.800 2309.710 1.000 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 818.750 -4.800 819.310 1.000 ;
    END
  END la_data_out[9]
  PIN la_oenb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 675.230 -4.800 675.790 1.000 ;
    END
  END la_oenb[0]
  PIN la_oenb[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2331.230 -4.800 2331.790 1.000 ;
    END
  END la_oenb[100]
  PIN la_oenb[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2347.790 -4.800 2348.350 1.000 ;
    END
  END la_oenb[101]
  PIN la_oenb[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2364.350 -4.800 2364.910 1.000 ;
    END
  END la_oenb[102]
  PIN la_oenb[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2380.910 -4.800 2381.470 1.000 ;
    END
  END la_oenb[103]
  PIN la_oenb[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2397.470 -4.800 2398.030 1.000 ;
    END
  END la_oenb[104]
  PIN la_oenb[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2414.030 -4.800 2414.590 1.000 ;
    END
  END la_oenb[105]
  PIN la_oenb[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2430.590 -4.800 2431.150 1.000 ;
    END
  END la_oenb[106]
  PIN la_oenb[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2447.150 -4.800 2447.710 1.000 ;
    END
  END la_oenb[107]
  PIN la_oenb[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2463.710 -4.800 2464.270 1.000 ;
    END
  END la_oenb[108]
  PIN la_oenb[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2480.270 -4.800 2480.830 1.000 ;
    END
  END la_oenb[109]
  PIN la_oenb[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 840.830 -4.800 841.390 1.000 ;
    END
  END la_oenb[10]
  PIN la_oenb[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2496.830 -4.800 2497.390 1.000 ;
    END
  END la_oenb[110]
  PIN la_oenb[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2513.390 -4.800 2513.950 1.000 ;
    END
  END la_oenb[111]
  PIN la_oenb[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2529.950 -4.800 2530.510 1.000 ;
    END
  END la_oenb[112]
  PIN la_oenb[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2546.510 -4.800 2547.070 1.000 ;
    END
  END la_oenb[113]
  PIN la_oenb[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2563.070 -4.800 2563.630 1.000 ;
    END
  END la_oenb[114]
  PIN la_oenb[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2579.630 -4.800 2580.190 1.000 ;
    END
  END la_oenb[115]
  PIN la_oenb[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2596.190 -4.800 2596.750 1.000 ;
    END
  END la_oenb[116]
  PIN la_oenb[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2612.750 -4.800 2613.310 1.000 ;
    END
  END la_oenb[117]
  PIN la_oenb[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2629.310 -4.800 2629.870 1.000 ;
    END
  END la_oenb[118]
  PIN la_oenb[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2645.870 -4.800 2646.430 1.000 ;
    END
  END la_oenb[119]
  PIN la_oenb[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 857.390 -4.800 857.950 1.000 ;
    END
  END la_oenb[11]
  PIN la_oenb[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2662.430 -4.800 2662.990 1.000 ;
    END
  END la_oenb[120]
  PIN la_oenb[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2678.990 -4.800 2679.550 1.000 ;
    END
  END la_oenb[121]
  PIN la_oenb[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2695.550 -4.800 2696.110 1.000 ;
    END
  END la_oenb[122]
  PIN la_oenb[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2712.110 -4.800 2712.670 1.000 ;
    END
  END la_oenb[123]
  PIN la_oenb[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2728.670 -4.800 2729.230 1.000 ;
    END
  END la_oenb[124]
  PIN la_oenb[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2745.230 -4.800 2745.790 1.000 ;
    END
  END la_oenb[125]
  PIN la_oenb[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2761.790 -4.800 2762.350 1.000 ;
    END
  END la_oenb[126]
  PIN la_oenb[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2778.350 -4.800 2778.910 1.000 ;
    END
  END la_oenb[127]
  PIN la_oenb[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 873.950 -4.800 874.510 1.000 ;
    END
  END la_oenb[12]
  PIN la_oenb[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 890.510 -4.800 891.070 1.000 ;
    END
  END la_oenb[13]
  PIN la_oenb[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 907.070 -4.800 907.630 1.000 ;
    END
  END la_oenb[14]
  PIN la_oenb[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 923.630 -4.800 924.190 1.000 ;
    END
  END la_oenb[15]
  PIN la_oenb[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 940.190 -4.800 940.750 1.000 ;
    END
  END la_oenb[16]
  PIN la_oenb[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 956.750 -4.800 957.310 1.000 ;
    END
  END la_oenb[17]
  PIN la_oenb[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 973.310 -4.800 973.870 1.000 ;
    END
  END la_oenb[18]
  PIN la_oenb[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 989.870 -4.800 990.430 1.000 ;
    END
  END la_oenb[19]
  PIN la_oenb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 691.790 -4.800 692.350 1.000 ;
    END
  END la_oenb[1]
  PIN la_oenb[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1006.430 -4.800 1006.990 1.000 ;
    END
  END la_oenb[20]
  PIN la_oenb[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1022.990 -4.800 1023.550 1.000 ;
    END
  END la_oenb[21]
  PIN la_oenb[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1039.550 -4.800 1040.110 1.000 ;
    END
  END la_oenb[22]
  PIN la_oenb[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1056.110 -4.800 1056.670 1.000 ;
    END
  END la_oenb[23]
  PIN la_oenb[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1072.670 -4.800 1073.230 1.000 ;
    END
  END la_oenb[24]
  PIN la_oenb[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1089.230 -4.800 1089.790 1.000 ;
    END
  END la_oenb[25]
  PIN la_oenb[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1105.790 -4.800 1106.350 1.000 ;
    END
  END la_oenb[26]
  PIN la_oenb[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1122.350 -4.800 1122.910 1.000 ;
    END
  END la_oenb[27]
  PIN la_oenb[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1138.910 -4.800 1139.470 1.000 ;
    END
  END la_oenb[28]
  PIN la_oenb[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1155.470 -4.800 1156.030 1.000 ;
    END
  END la_oenb[29]
  PIN la_oenb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 708.350 -4.800 708.910 1.000 ;
    END
  END la_oenb[2]
  PIN la_oenb[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1172.030 -4.800 1172.590 1.000 ;
    END
  END la_oenb[30]
  PIN la_oenb[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1188.590 -4.800 1189.150 1.000 ;
    END
  END la_oenb[31]
  PIN la_oenb[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1205.150 -4.800 1205.710 1.000 ;
    END
  END la_oenb[32]
  PIN la_oenb[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1221.710 -4.800 1222.270 1.000 ;
    END
  END la_oenb[33]
  PIN la_oenb[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1238.270 -4.800 1238.830 1.000 ;
    END
  END la_oenb[34]
  PIN la_oenb[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1254.830 -4.800 1255.390 1.000 ;
    END
  END la_oenb[35]
  PIN la_oenb[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1271.390 -4.800 1271.950 1.000 ;
    END
  END la_oenb[36]
  PIN la_oenb[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1287.950 -4.800 1288.510 1.000 ;
    END
  END la_oenb[37]
  PIN la_oenb[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1304.510 -4.800 1305.070 1.000 ;
    END
  END la_oenb[38]
  PIN la_oenb[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1321.070 -4.800 1321.630 1.000 ;
    END
  END la_oenb[39]
  PIN la_oenb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 724.910 -4.800 725.470 1.000 ;
    END
  END la_oenb[3]
  PIN la_oenb[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1337.630 -4.800 1338.190 1.000 ;
    END
  END la_oenb[40]
  PIN la_oenb[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1354.190 -4.800 1354.750 1.000 ;
    END
  END la_oenb[41]
  PIN la_oenb[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1370.750 -4.800 1371.310 1.000 ;
    END
  END la_oenb[42]
  PIN la_oenb[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1387.310 -4.800 1387.870 1.000 ;
    END
  END la_oenb[43]
  PIN la_oenb[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1403.870 -4.800 1404.430 1.000 ;
    END
  END la_oenb[44]
  PIN la_oenb[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1420.430 -4.800 1420.990 1.000 ;
    END
  END la_oenb[45]
  PIN la_oenb[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1436.990 -4.800 1437.550 1.000 ;
    END
  END la_oenb[46]
  PIN la_oenb[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1453.550 -4.800 1454.110 1.000 ;
    END
  END la_oenb[47]
  PIN la_oenb[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1470.110 -4.800 1470.670 1.000 ;
    END
  END la_oenb[48]
  PIN la_oenb[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1486.670 -4.800 1487.230 1.000 ;
    END
  END la_oenb[49]
  PIN la_oenb[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 741.470 -4.800 742.030 1.000 ;
    END
  END la_oenb[4]
  PIN la_oenb[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1503.230 -4.800 1503.790 1.000 ;
    END
  END la_oenb[50]
  PIN la_oenb[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1519.790 -4.800 1520.350 1.000 ;
    END
  END la_oenb[51]
  PIN la_oenb[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1536.350 -4.800 1536.910 1.000 ;
    END
  END la_oenb[52]
  PIN la_oenb[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1552.910 -4.800 1553.470 1.000 ;
    END
  END la_oenb[53]
  PIN la_oenb[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1569.470 -4.800 1570.030 1.000 ;
    END
  END la_oenb[54]
  PIN la_oenb[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1586.030 -4.800 1586.590 1.000 ;
    END
  END la_oenb[55]
  PIN la_oenb[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1602.590 -4.800 1603.150 1.000 ;
    END
  END la_oenb[56]
  PIN la_oenb[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1619.150 -4.800 1619.710 1.000 ;
    END
  END la_oenb[57]
  PIN la_oenb[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1635.710 -4.800 1636.270 1.000 ;
    END
  END la_oenb[58]
  PIN la_oenb[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1652.270 -4.800 1652.830 1.000 ;
    END
  END la_oenb[59]
  PIN la_oenb[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 758.030 -4.800 758.590 1.000 ;
    END
  END la_oenb[5]
  PIN la_oenb[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1668.830 -4.800 1669.390 1.000 ;
    END
  END la_oenb[60]
  PIN la_oenb[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1685.390 -4.800 1685.950 1.000 ;
    END
  END la_oenb[61]
  PIN la_oenb[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1701.950 -4.800 1702.510 1.000 ;
    END
  END la_oenb[62]
  PIN la_oenb[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1718.510 -4.800 1719.070 1.000 ;
    END
  END la_oenb[63]
  PIN la_oenb[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1735.070 -4.800 1735.630 1.000 ;
    END
  END la_oenb[64]
  PIN la_oenb[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1751.630 -4.800 1752.190 1.000 ;
    END
  END la_oenb[65]
  PIN la_oenb[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1768.190 -4.800 1768.750 1.000 ;
    END
  END la_oenb[66]
  PIN la_oenb[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1784.750 -4.800 1785.310 1.000 ;
    END
  END la_oenb[67]
  PIN la_oenb[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1801.310 -4.800 1801.870 1.000 ;
    END
  END la_oenb[68]
  PIN la_oenb[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1817.870 -4.800 1818.430 1.000 ;
    END
  END la_oenb[69]
  PIN la_oenb[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 774.590 -4.800 775.150 1.000 ;
    END
  END la_oenb[6]
  PIN la_oenb[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1834.430 -4.800 1834.990 1.000 ;
    END
  END la_oenb[70]
  PIN la_oenb[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1850.990 -4.800 1851.550 1.000 ;
    END
  END la_oenb[71]
  PIN la_oenb[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1867.550 -4.800 1868.110 1.000 ;
    END
  END la_oenb[72]
  PIN la_oenb[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1884.110 -4.800 1884.670 1.000 ;
    END
  END la_oenb[73]
  PIN la_oenb[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1900.670 -4.800 1901.230 1.000 ;
    END
  END la_oenb[74]
  PIN la_oenb[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1917.230 -4.800 1917.790 1.000 ;
    END
  END la_oenb[75]
  PIN la_oenb[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1933.790 -4.800 1934.350 1.000 ;
    END
  END la_oenb[76]
  PIN la_oenb[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1950.350 -4.800 1950.910 1.000 ;
    END
  END la_oenb[77]
  PIN la_oenb[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1966.910 -4.800 1967.470 1.000 ;
    END
  END la_oenb[78]
  PIN la_oenb[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1983.470 -4.800 1984.030 1.000 ;
    END
  END la_oenb[79]
  PIN la_oenb[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 791.150 -4.800 791.710 1.000 ;
    END
  END la_oenb[7]
  PIN la_oenb[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2000.030 -4.800 2000.590 1.000 ;
    END
  END la_oenb[80]
  PIN la_oenb[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2016.590 -4.800 2017.150 1.000 ;
    END
  END la_oenb[81]
  PIN la_oenb[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2033.150 -4.800 2033.710 1.000 ;
    END
  END la_oenb[82]
  PIN la_oenb[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2049.710 -4.800 2050.270 1.000 ;
    END
  END la_oenb[83]
  PIN la_oenb[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2066.270 -4.800 2066.830 1.000 ;
    END
  END la_oenb[84]
  PIN la_oenb[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2082.830 -4.800 2083.390 1.000 ;
    END
  END la_oenb[85]
  PIN la_oenb[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2099.390 -4.800 2099.950 1.000 ;
    END
  END la_oenb[86]
  PIN la_oenb[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2115.950 -4.800 2116.510 1.000 ;
    END
  END la_oenb[87]
  PIN la_oenb[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2132.510 -4.800 2133.070 1.000 ;
    END
  END la_oenb[88]
  PIN la_oenb[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2149.070 -4.800 2149.630 1.000 ;
    END
  END la_oenb[89]
  PIN la_oenb[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 807.710 -4.800 808.270 1.000 ;
    END
  END la_oenb[8]
  PIN la_oenb[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2165.630 -4.800 2166.190 1.000 ;
    END
  END la_oenb[90]
  PIN la_oenb[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2182.190 -4.800 2182.750 1.000 ;
    END
  END la_oenb[91]
  PIN la_oenb[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2198.750 -4.800 2199.310 1.000 ;
    END
  END la_oenb[92]
  PIN la_oenb[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2215.310 -4.800 2215.870 1.000 ;
    END
  END la_oenb[93]
  PIN la_oenb[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2231.870 -4.800 2232.430 1.000 ;
    END
  END la_oenb[94]
  PIN la_oenb[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2248.430 -4.800 2248.990 1.000 ;
    END
  END la_oenb[95]
  PIN la_oenb[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2264.990 -4.800 2265.550 1.000 ;
    END
  END la_oenb[96]
  PIN la_oenb[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2281.550 -4.800 2282.110 1.000 ;
    END
  END la_oenb[97]
  PIN la_oenb[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2298.110 -4.800 2298.670 1.000 ;
    END
  END la_oenb[98]
  PIN la_oenb[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2314.670 -4.800 2315.230 1.000 ;
    END
  END la_oenb[99]
  PIN la_oenb[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 824.270 -4.800 824.830 1.000 ;
    END
  END la_oenb[9]
  PIN user_clock2
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2783.870 -4.800 2784.430 1.000 ;
    END
  END user_clock2
  PIN user_irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2789.390 -4.800 2789.950 1.000 ;
    END
  END user_irq[0]
  PIN user_irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2794.910 -4.800 2795.470 1.000 ;
    END
  END user_irq[1]
  PIN user_irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2800.430 -4.800 2800.990 1.000 ;
    END
  END user_irq[2]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 8.970 10.640 12.070 3468.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 188.970 10.640 192.070 115.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 188.970 551.540 192.070 680.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 188.970 1116.540 192.070 1260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 188.970 1696.540 192.070 1820.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 188.970 2256.540 192.070 2415.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 188.970 2851.540 192.070 2975.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 188.970 3411.540 192.070 3468.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 368.970 10.640 372.070 115.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 368.970 551.540 372.070 680.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 368.970 1116.540 372.070 1260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 368.970 1696.540 372.070 1820.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 368.970 2256.540 372.070 2415.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 368.970 2851.540 372.070 2975.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 368.970 3411.540 372.070 3468.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 548.970 10.640 552.070 115.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 548.970 551.540 552.070 680.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 548.970 1116.540 552.070 1260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 548.970 1696.540 552.070 1820.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 548.970 2256.540 552.070 2415.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 548.970 2851.540 552.070 2975.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 548.970 3411.540 552.070 3468.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 728.970 10.640 732.070 115.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 728.970 551.540 732.070 680.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 728.970 1116.540 732.070 1260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 728.970 1696.540 732.070 1820.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 728.970 2256.540 732.070 2415.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 728.970 2851.540 732.070 2975.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 728.970 3411.540 732.070 3468.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 908.970 10.640 912.070 140.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 908.970 557.500 912.070 2940.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 908.970 3357.500 912.070 3468.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 1088.970 10.640 1092.070 140.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1088.970 557.500 1092.070 2940.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1088.970 3357.500 1092.070 3468.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 1268.970 10.640 1272.070 140.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1268.970 557.500 1272.070 2940.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1268.970 3357.500 1272.070 3468.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 1448.970 10.640 1452.070 3468.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 1628.970 10.640 1632.070 140.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1628.970 557.500 1632.070 2940.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1628.970 3357.500 1632.070 3468.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 1808.970 10.640 1812.070 140.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1808.970 557.500 1812.070 2940.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1808.970 3357.500 1812.070 3468.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 1988.970 10.640 1992.070 3468.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 2168.970 10.640 2172.070 115.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2168.970 551.540 2172.070 680.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2168.970 1116.540 2172.070 1260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2168.970 1696.540 2172.070 1820.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2168.970 2256.540 2172.070 2415.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2168.970 2851.540 2172.070 2975.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2168.970 3411.540 2172.070 3468.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 2348.970 10.640 2352.070 115.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2348.970 551.540 2352.070 680.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2348.970 1116.540 2352.070 1260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2348.970 1696.540 2352.070 1820.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2348.970 2256.540 2352.070 2415.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2348.970 2851.540 2352.070 2975.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2348.970 3411.540 2352.070 3468.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 2528.970 10.640 2532.070 115.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2528.970 551.540 2532.070 680.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2528.970 1116.540 2532.070 1260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2528.970 1696.540 2532.070 1820.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2528.970 2256.540 2532.070 2415.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2528.970 2851.540 2532.070 2975.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2528.970 3411.540 2532.070 3468.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 2708.970 10.640 2712.070 115.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2708.970 551.540 2712.070 680.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2708.970 1116.540 2712.070 1260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2708.970 1696.540 2712.070 1820.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2708.970 2256.540 2712.070 2415.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2708.970 2851.540 2712.070 2975.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2708.970 3411.540 2712.070 3468.240 ;
    END
#    PORT
#      LAYER met5 ;
#        RECT 5.280 14.330 2874.320 17.430 ;
#    END
#    PORT
#      LAYER met5 ;
#        RECT 5.280 194.330 2874.320 197.430 ;
#    END
#    PORT
#      LAYER met5 ;
#        RECT 5.280 374.330 2874.320 377.430 ;
#    END
#    PORT
#      LAYER met5 ;
#        RECT 5.280 554.330 2874.320 557.430 ;
#    END
#    PORT
#      LAYER met5 ;
#        RECT 5.280 734.330 2874.320 737.430 ;
#    END
#    PORT
#      LAYER met5 ;
#        RECT 5.280 914.330 2874.320 917.430 ;
#    END
#    PORT
#      LAYER met5 ;
#        RECT 5.280 1094.330 2874.320 1097.430 ;
#    END
#    PORT
#      LAYER met5 ;
#        RECT 5.280 1274.330 2874.320 1277.430 ;
#    END
#    PORT
#      LAYER met5 ;
#        RECT 5.280 1454.330 2874.320 1457.430 ;
#    END
#    PORT
#      LAYER met5 ;
#        RECT 5.280 1634.330 2874.320 1637.430 ;
#    END
#    PORT
#      LAYER met5 ;
#        RECT 5.280 1814.330 2874.320 1817.430 ;
#    END
#    PORT
#      LAYER met5 ;
#        RECT 5.280 1994.330 2874.320 1997.430 ;
#    END
#    PORT
#      LAYER met5 ;
#        RECT 5.280 2174.330 2874.320 2177.430 ;
#    END
#    PORT
#      LAYER met5 ;
#        RECT 5.280 2354.330 2874.320 2357.430 ;
#    END
#    PORT
#      LAYER met5 ;
#        RECT 5.280 2534.330 2874.320 2537.430 ;
#    END
#    PORT
#      LAYER met5 ;
#        RECT 5.280 2714.330 2874.320 2717.430 ;
#    END
#    PORT
#      LAYER met5 ;
#        RECT 5.280 2894.330 2874.320 2897.430 ;
#    END
#    PORT
#      LAYER met5 ;
#        RECT 5.280 3074.330 2874.320 3077.430 ;
#    END
#    PORT
#      LAYER met5 ;
#        RECT 5.280 3254.330 2874.320 3257.430 ;
#    END
#    PORT
#      LAYER met5 ;
#        RECT 5.280 3434.330 2874.320 3437.430 ;
#    END
    PORT
      LAYER met4 ;
        RECT 845.310 2972.720 848.410 3359.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 2831.590 677.040 2834.690 1118.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 845.310 138.480 848.410 552.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 2831.590 1259.120 2834.690 1700.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 2831.590 1819.440 2834.690 2260.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 2831.590 111.280 2834.690 552.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 2831.590 2972.720 2834.690 3413.840 ;
    END
    PORT
      LAYER met4 ;
        RECT 2831.590 2412.400 2834.690 2853.520 ;
    END
#    PORT
#      LAYER met5 ;
#        RECT 1988.970 1149.350 2874.320 1152.450 ;
#    END
#    PORT
#      LAYER met5 ;
#        RECT 8.970 1149.350 912.070 1152.450 ;
#    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 98.970 10.640 102.070 115.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 98.970 551.540 102.070 680.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 98.970 1116.540 102.070 1260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 98.970 1696.540 102.070 1820.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 98.970 2256.540 102.070 2415.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 98.970 2851.540 102.070 2975.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 98.970 3411.540 102.070 3468.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 278.970 10.640 282.070 115.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 278.970 551.540 282.070 680.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 278.970 1116.540 282.070 1260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 278.970 1696.540 282.070 1820.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 278.970 2256.540 282.070 2415.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 278.970 2851.540 282.070 2975.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 278.970 3411.540 282.070 3468.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 458.970 10.640 462.070 115.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 458.970 551.540 462.070 680.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 458.970 1116.540 462.070 1260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 458.970 1696.540 462.070 1820.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 458.970 2256.540 462.070 2415.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 458.970 2851.540 462.070 2975.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 458.970 3411.540 462.070 3468.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 638.970 10.640 642.070 115.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 638.970 551.540 642.070 680.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 638.970 1116.540 642.070 1260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 638.970 1696.540 642.070 1820.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 638.970 2256.540 642.070 2415.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 638.970 2851.540 642.070 2975.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 638.970 3411.540 642.070 3468.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 818.970 10.640 822.070 3468.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 998.970 10.640 1002.070 140.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 998.970 557.500 1002.070 2940.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 998.970 3357.500 1002.070 3468.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 1178.970 10.640 1182.070 140.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1178.970 557.500 1182.070 2940.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1178.970 3357.500 1182.070 3468.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 1358.970 10.640 1362.070 140.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1358.970 557.500 1362.070 2940.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1358.970 3357.500 1362.070 3468.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 1538.970 10.640 1542.070 140.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1538.970 557.500 1542.070 2940.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1538.970 3357.500 1542.070 3468.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 1718.970 10.640 1722.070 140.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1718.970 557.500 1722.070 2940.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1718.970 3357.500 1722.070 3468.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 1898.970 10.640 1902.070 140.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1898.970 557.500 1902.070 2940.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 1898.970 3357.500 1902.070 3468.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 2078.970 10.640 2082.070 3468.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 2258.970 10.640 2262.070 115.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2258.970 551.540 2262.070 680.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2258.970 1116.540 2262.070 1260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2258.970 1696.540 2262.070 1820.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2258.970 2256.540 2262.070 2415.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2258.970 2851.540 2262.070 2975.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2258.970 3411.540 2262.070 3468.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 2438.970 10.640 2442.070 115.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2438.970 551.540 2442.070 680.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2438.970 1116.540 2442.070 1260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2438.970 1696.540 2442.070 1820.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2438.970 2256.540 2442.070 2415.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2438.970 2851.540 2442.070 2975.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2438.970 3411.540 2442.070 3468.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 2618.970 10.640 2622.070 115.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2618.970 551.540 2622.070 680.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2618.970 1116.540 2622.070 1260.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2618.970 1696.540 2622.070 1820.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2618.970 2256.540 2622.070 2415.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2618.970 2851.540 2622.070 2975.000 ;
    END
    PORT
      LAYER met4 ;
        RECT 2618.970 3411.540 2622.070 3468.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 2798.970 10.640 2802.070 3468.240 ;
    END
#    PORT
#      LAYER met5 ;
#        RECT 5.280 104.330 2874.320 107.430 ;
#    END
#    PORT
#      LAYER met5 ;
#        RECT 5.280 284.330 2874.320 287.430 ;
#    END
#    PORT
#      LAYER met5 ;
#        RECT 5.280 464.330 2874.320 467.430 ;
#    END
#    PORT
#      LAYER met5 ;
#        RECT 5.280 644.330 2874.320 647.430 ;
#    END
#    PORT
#      LAYER met5 ;
#        RECT 5.280 824.330 2874.320 827.430 ;
#    END
#    PORT
#      LAYER met5 ;
#        RECT 5.280 1004.330 2874.320 1007.430 ;
#    END
#    PORT
#      LAYER met5 ;
#        RECT 5.280 1184.330 2874.320 1187.430 ;
#    END
#    PORT
#      LAYER met5 ;
#        RECT 5.280 1364.330 2874.320 1367.430 ;
#    END
#    PORT
#      LAYER met5 ;
#        RECT 5.280 1544.330 2874.320 1547.430 ;
#    END
#    PORT
#      LAYER met5 ;
#        RECT 5.280 1724.330 2874.320 1727.430 ;
#    END
#    PORT
#      LAYER met5 ;
#        RECT 5.280 1904.330 2874.320 1907.430 ;
#    END
#    PORT
#      LAYER met5 ;
#        RECT 5.280 2084.330 2874.320 2087.430 ;
#    END
#    PORT
#      LAYER met5 ;
#        RECT 5.280 2264.330 2874.320 2267.430 ;
#    END
#    PORT
#      LAYER met5 ;
#        RECT 5.280 2444.330 2874.320 2447.430 ;
#    END
#    PORT
#      LAYER met5 ;
#        RECT 5.280 2624.330 2874.320 2627.430 ;
#    END
#    PORT
#      LAYER met5 ;
#        RECT 5.280 2804.330 2874.320 2807.430 ;
#    END
#    PORT
#      LAYER met5 ;
#        RECT 5.280 2984.330 2874.320 2987.430 ;
#    END
#    PORT
#      LAYER met5 ;
#        RECT 5.280 3164.330 2874.320 3167.430 ;
#    END
#    PORT
#      LAYER met5 ;
#        RECT 5.280 3344.330 2874.320 3347.430 ;
#    END
    PORT
      LAYER met4 ;
        RECT 45.830 114.000 48.930 555.120 ;
    END
    PORT
      LAYER met4 ;
        RECT 45.830 679.760 48.930 1120.880 ;
    END
    PORT
      LAYER met4 ;
        RECT 1437.790 2937.360 1440.890 3362.160 ;
    END
    PORT
      LAYER met4 ;
        RECT 45.830 1256.400 48.930 1697.520 ;
    END
    PORT
      LAYER met4 ;
        RECT 1437.790 135.760 1440.890 560.560 ;
    END
    PORT
      LAYER met4 ;
        RECT 45.830 1816.720 48.930 2257.840 ;
    END
#    PORT
#      LAYER met5 ;
#        RECT 818.970 3410.350 2082.070 3413.450 ;
#    END
    PORT
      LAYER met4 ;
        RECT 45.830 2409.680 48.930 2856.240 ;
    END
    PORT
      LAYER met4 ;
        RECT 45.830 2970.000 48.930 3416.560 ;
    END
#    PORT
#      LAYER met5 ;
#        RECT 5.280 2910.550 822.070 2913.650 ;
#    END
#    PORT
#      LAYER met5 ;
#        RECT 5.280 3423.950 822.070 3427.050 ;
#    END
#    PORT
#      LAYER met5 ;
#        RECT 2078.970 2910.550 2802.070 2913.650 ;
#    END
#    PORT
#      LAYER met5 ;
#        RECT 2078.970 3423.950 2802.070 3427.050 ;
#    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 79.070 -4.800 79.630 1.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 84.590 -4.800 85.150 1.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.110 -4.800 90.670 1.000 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.190 -4.800 112.750 1.000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.870 -4.800 300.430 1.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 316.430 -4.800 316.990 1.000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 332.990 -4.800 333.550 1.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 349.550 -4.800 350.110 1.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 366.110 -4.800 366.670 1.000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 382.670 -4.800 383.230 1.000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 399.230 -4.800 399.790 1.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 415.790 -4.800 416.350 1.000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 432.350 -4.800 432.910 1.000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 448.910 -4.800 449.470 1.000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 134.270 -4.800 134.830 1.000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 465.470 -4.800 466.030 1.000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 482.030 -4.800 482.590 1.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 498.590 -4.800 499.150 1.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 515.150 -4.800 515.710 1.000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 531.710 -4.800 532.270 1.000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 548.270 -4.800 548.830 1.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 564.830 -4.800 565.390 1.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 581.390 -4.800 581.950 1.000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 597.950 -4.800 598.510 1.000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 614.510 -4.800 615.070 1.000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.350 -4.800 156.910 1.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 631.070 -4.800 631.630 1.000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 647.630 -4.800 648.190 1.000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 178.430 -4.800 178.990 1.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 200.510 -4.800 201.070 1.000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 217.070 -4.800 217.630 1.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.630 -4.800 234.190 1.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 250.190 -4.800 250.750 1.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 266.750 -4.800 267.310 1.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.310 -4.800 283.870 1.000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 95.630 -4.800 96.190 1.000 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 117.710 -4.800 118.270 1.000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.390 -4.800 305.950 1.000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 321.950 -4.800 322.510 1.000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 338.510 -4.800 339.070 1.000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 355.070 -4.800 355.630 1.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 371.630 -4.800 372.190 1.000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 388.190 -4.800 388.750 1.000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 404.750 -4.800 405.310 1.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 421.310 -4.800 421.870 1.000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 437.870 -4.800 438.430 1.000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 454.430 -4.800 454.990 1.000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.790 -4.800 140.350 1.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 470.990 -4.800 471.550 1.000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 487.550 -4.800 488.110 1.000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 504.110 -4.800 504.670 1.000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 520.670 -4.800 521.230 1.000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 537.230 -4.800 537.790 1.000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 553.790 -4.800 554.350 1.000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 570.350 -4.800 570.910 1.000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 586.910 -4.800 587.470 1.000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 603.470 -4.800 604.030 1.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 620.030 -4.800 620.590 1.000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.870 -4.800 162.430 1.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 636.590 -4.800 637.150 1.000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 653.150 -4.800 653.710 1.000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.950 -4.800 184.510 1.000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 206.030 -4.800 206.590 1.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.590 -4.800 223.150 1.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 239.150 -4.800 239.710 1.000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 255.710 -4.800 256.270 1.000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 272.270 -4.800 272.830 1.000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.830 -4.800 289.390 1.000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 123.230 -4.800 123.790 1.000 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 310.910 -4.800 311.470 1.000 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 327.470 -4.800 328.030 1.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 344.030 -4.800 344.590 1.000 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 360.590 -4.800 361.150 1.000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 377.150 -4.800 377.710 1.000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 393.710 -4.800 394.270 1.000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 410.270 -4.800 410.830 1.000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 426.830 -4.800 427.390 1.000 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 443.390 -4.800 443.950 1.000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 459.950 -4.800 460.510 1.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 145.310 -4.800 145.870 1.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 476.510 -4.800 477.070 1.000 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 493.070 -4.800 493.630 1.000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 509.630 -4.800 510.190 1.000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 526.190 -4.800 526.750 1.000 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 542.750 -4.800 543.310 1.000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 559.310 -4.800 559.870 1.000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 575.870 -4.800 576.430 1.000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 592.430 -4.800 592.990 1.000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 608.990 -4.800 609.550 1.000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 625.550 -4.800 626.110 1.000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.390 -4.800 167.950 1.000 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 642.110 -4.800 642.670 1.000 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 658.670 -4.800 659.230 1.000 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 189.470 -4.800 190.030 1.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 211.550 -4.800 212.110 1.000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.110 -4.800 228.670 1.000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.670 -4.800 245.230 1.000 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 261.230 -4.800 261.790 1.000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 277.790 -4.800 278.350 1.000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.350 -4.800 294.910 1.000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.750 -4.800 129.310 1.000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.830 -4.800 151.390 1.000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 172.910 -4.800 173.470 1.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 194.990 -4.800 195.550 1.000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.150 -4.800 101.710 1.000 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.670 -4.800 107.230 1.000 ;
    END
  END wbs_we_i
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 2874.080 3468.085 ;
      LAYER met1 ;
        RECT 5.520 6.840 2874.080 3468.240 ;
      LAYER met2 ;
        RECT 6.990 3478.720 46.590 3479.000 ;
        RECT 47.710 3478.720 126.170 3479.000 ;
        RECT 127.290 3478.720 205.750 3479.000 ;
        RECT 206.870 3478.720 285.330 3479.000 ;
        RECT 286.450 3478.720 364.910 3479.000 ;
        RECT 366.030 3478.720 444.490 3479.000 ;
        RECT 445.610 3478.720 524.070 3479.000 ;
        RECT 525.190 3478.720 603.650 3479.000 ;
        RECT 604.770 3478.720 683.230 3479.000 ;
        RECT 684.350 3478.720 762.810 3479.000 ;
        RECT 763.930 3478.720 842.390 3479.000 ;
        RECT 843.510 3478.720 921.970 3479.000 ;
        RECT 923.090 3478.720 1001.550 3479.000 ;
        RECT 1002.670 3478.720 1081.130 3479.000 ;
        RECT 1082.250 3478.720 1160.710 3479.000 ;
        RECT 1161.830 3478.720 1240.290 3479.000 ;
        RECT 1241.410 3478.720 1319.870 3479.000 ;
        RECT 1320.990 3478.720 1399.450 3479.000 ;
        RECT 1400.570 3478.720 1479.030 3479.000 ;
        RECT 1480.150 3478.720 1558.610 3479.000 ;
        RECT 1559.730 3478.720 1638.190 3479.000 ;
        RECT 1639.310 3478.720 1717.770 3479.000 ;
        RECT 1718.890 3478.720 1797.350 3479.000 ;
        RECT 1798.470 3478.720 1876.930 3479.000 ;
        RECT 1878.050 3478.720 1956.510 3479.000 ;
        RECT 1957.630 3478.720 2036.090 3479.000 ;
        RECT 2037.210 3478.720 2115.670 3479.000 ;
        RECT 2116.790 3478.720 2195.250 3479.000 ;
        RECT 2196.370 3478.720 2274.830 3479.000 ;
        RECT 2275.950 3478.720 2354.410 3479.000 ;
        RECT 2355.530 3478.720 2433.990 3479.000 ;
        RECT 2435.110 3478.720 2513.570 3479.000 ;
        RECT 2514.690 3478.720 2593.150 3479.000 ;
        RECT 2594.270 3478.720 2672.730 3479.000 ;
        RECT 2673.850 3478.720 2752.310 3479.000 ;
        RECT 2753.430 3478.720 2831.890 3479.000 ;
        RECT 2833.010 3478.720 2871.690 3479.000 ;
        RECT 6.990 1.280 2871.690 3478.720 ;
        RECT 6.990 0.270 78.790 1.280 ;
        RECT 79.910 0.270 84.310 1.280 ;
        RECT 85.430 0.270 89.830 1.280 ;
        RECT 90.950 0.270 95.350 1.280 ;
        RECT 96.470 0.270 100.870 1.280 ;
        RECT 101.990 0.270 106.390 1.280 ;
        RECT 107.510 0.270 111.910 1.280 ;
        RECT 113.030 0.270 117.430 1.280 ;
        RECT 118.550 0.270 122.950 1.280 ;
        RECT 124.070 0.270 128.470 1.280 ;
        RECT 129.590 0.270 133.990 1.280 ;
        RECT 135.110 0.270 139.510 1.280 ;
        RECT 140.630 0.270 145.030 1.280 ;
        RECT 146.150 0.270 150.550 1.280 ;
        RECT 151.670 0.270 156.070 1.280 ;
        RECT 157.190 0.270 161.590 1.280 ;
        RECT 162.710 0.270 167.110 1.280 ;
        RECT 168.230 0.270 172.630 1.280 ;
        RECT 173.750 0.270 178.150 1.280 ;
        RECT 179.270 0.270 183.670 1.280 ;
        RECT 184.790 0.270 189.190 1.280 ;
        RECT 190.310 0.270 194.710 1.280 ;
        RECT 195.830 0.270 200.230 1.280 ;
        RECT 201.350 0.270 205.750 1.280 ;
        RECT 206.870 0.270 211.270 1.280 ;
        RECT 212.390 0.270 216.790 1.280 ;
        RECT 217.910 0.270 222.310 1.280 ;
        RECT 223.430 0.270 227.830 1.280 ;
        RECT 228.950 0.270 233.350 1.280 ;
        RECT 234.470 0.270 238.870 1.280 ;
        RECT 239.990 0.270 244.390 1.280 ;
        RECT 245.510 0.270 249.910 1.280 ;
        RECT 251.030 0.270 255.430 1.280 ;
        RECT 256.550 0.270 260.950 1.280 ;
        RECT 262.070 0.270 266.470 1.280 ;
        RECT 267.590 0.270 271.990 1.280 ;
        RECT 273.110 0.270 277.510 1.280 ;
        RECT 278.630 0.270 283.030 1.280 ;
        RECT 284.150 0.270 288.550 1.280 ;
        RECT 289.670 0.270 294.070 1.280 ;
        RECT 295.190 0.270 299.590 1.280 ;
        RECT 300.710 0.270 305.110 1.280 ;
        RECT 306.230 0.270 310.630 1.280 ;
        RECT 311.750 0.270 316.150 1.280 ;
        RECT 317.270 0.270 321.670 1.280 ;
        RECT 322.790 0.270 327.190 1.280 ;
        RECT 328.310 0.270 332.710 1.280 ;
        RECT 333.830 0.270 338.230 1.280 ;
        RECT 339.350 0.270 343.750 1.280 ;
        RECT 344.870 0.270 349.270 1.280 ;
        RECT 350.390 0.270 354.790 1.280 ;
        RECT 355.910 0.270 360.310 1.280 ;
        RECT 361.430 0.270 365.830 1.280 ;
        RECT 366.950 0.270 371.350 1.280 ;
        RECT 372.470 0.270 376.870 1.280 ;
        RECT 377.990 0.270 382.390 1.280 ;
        RECT 383.510 0.270 387.910 1.280 ;
        RECT 389.030 0.270 393.430 1.280 ;
        RECT 394.550 0.270 398.950 1.280 ;
        RECT 400.070 0.270 404.470 1.280 ;
        RECT 405.590 0.270 409.990 1.280 ;
        RECT 411.110 0.270 415.510 1.280 ;
        RECT 416.630 0.270 421.030 1.280 ;
        RECT 422.150 0.270 426.550 1.280 ;
        RECT 427.670 0.270 432.070 1.280 ;
        RECT 433.190 0.270 437.590 1.280 ;
        RECT 438.710 0.270 443.110 1.280 ;
        RECT 444.230 0.270 448.630 1.280 ;
        RECT 449.750 0.270 454.150 1.280 ;
        RECT 455.270 0.270 459.670 1.280 ;
        RECT 460.790 0.270 465.190 1.280 ;
        RECT 466.310 0.270 470.710 1.280 ;
        RECT 471.830 0.270 476.230 1.280 ;
        RECT 477.350 0.270 481.750 1.280 ;
        RECT 482.870 0.270 487.270 1.280 ;
        RECT 488.390 0.270 492.790 1.280 ;
        RECT 493.910 0.270 498.310 1.280 ;
        RECT 499.430 0.270 503.830 1.280 ;
        RECT 504.950 0.270 509.350 1.280 ;
        RECT 510.470 0.270 514.870 1.280 ;
        RECT 515.990 0.270 520.390 1.280 ;
        RECT 521.510 0.270 525.910 1.280 ;
        RECT 527.030 0.270 531.430 1.280 ;
        RECT 532.550 0.270 536.950 1.280 ;
        RECT 538.070 0.270 542.470 1.280 ;
        RECT 543.590 0.270 547.990 1.280 ;
        RECT 549.110 0.270 553.510 1.280 ;
        RECT 554.630 0.270 559.030 1.280 ;
        RECT 560.150 0.270 564.550 1.280 ;
        RECT 565.670 0.270 570.070 1.280 ;
        RECT 571.190 0.270 575.590 1.280 ;
        RECT 576.710 0.270 581.110 1.280 ;
        RECT 582.230 0.270 586.630 1.280 ;
        RECT 587.750 0.270 592.150 1.280 ;
        RECT 593.270 0.270 597.670 1.280 ;
        RECT 598.790 0.270 603.190 1.280 ;
        RECT 604.310 0.270 608.710 1.280 ;
        RECT 609.830 0.270 614.230 1.280 ;
        RECT 615.350 0.270 619.750 1.280 ;
        RECT 620.870 0.270 625.270 1.280 ;
        RECT 626.390 0.270 630.790 1.280 ;
        RECT 631.910 0.270 636.310 1.280 ;
        RECT 637.430 0.270 641.830 1.280 ;
        RECT 642.950 0.270 647.350 1.280 ;
        RECT 648.470 0.270 652.870 1.280 ;
        RECT 653.990 0.270 658.390 1.280 ;
        RECT 659.510 0.270 663.910 1.280 ;
        RECT 665.030 0.270 669.430 1.280 ;
        RECT 670.550 0.270 674.950 1.280 ;
        RECT 676.070 0.270 680.470 1.280 ;
        RECT 681.590 0.270 685.990 1.280 ;
        RECT 687.110 0.270 691.510 1.280 ;
        RECT 692.630 0.270 697.030 1.280 ;
        RECT 698.150 0.270 702.550 1.280 ;
        RECT 703.670 0.270 708.070 1.280 ;
        RECT 709.190 0.270 713.590 1.280 ;
        RECT 714.710 0.270 719.110 1.280 ;
        RECT 720.230 0.270 724.630 1.280 ;
        RECT 725.750 0.270 730.150 1.280 ;
        RECT 731.270 0.270 735.670 1.280 ;
        RECT 736.790 0.270 741.190 1.280 ;
        RECT 742.310 0.270 746.710 1.280 ;
        RECT 747.830 0.270 752.230 1.280 ;
        RECT 753.350 0.270 757.750 1.280 ;
        RECT 758.870 0.270 763.270 1.280 ;
        RECT 764.390 0.270 768.790 1.280 ;
        RECT 769.910 0.270 774.310 1.280 ;
        RECT 775.430 0.270 779.830 1.280 ;
        RECT 780.950 0.270 785.350 1.280 ;
        RECT 786.470 0.270 790.870 1.280 ;
        RECT 791.990 0.270 796.390 1.280 ;
        RECT 797.510 0.270 801.910 1.280 ;
        RECT 803.030 0.270 807.430 1.280 ;
        RECT 808.550 0.270 812.950 1.280 ;
        RECT 814.070 0.270 818.470 1.280 ;
        RECT 819.590 0.270 823.990 1.280 ;
        RECT 825.110 0.270 829.510 1.280 ;
        RECT 830.630 0.270 835.030 1.280 ;
        RECT 836.150 0.270 840.550 1.280 ;
        RECT 841.670 0.270 846.070 1.280 ;
        RECT 847.190 0.270 851.590 1.280 ;
        RECT 852.710 0.270 857.110 1.280 ;
        RECT 858.230 0.270 862.630 1.280 ;
        RECT 863.750 0.270 868.150 1.280 ;
        RECT 869.270 0.270 873.670 1.280 ;
        RECT 874.790 0.270 879.190 1.280 ;
        RECT 880.310 0.270 884.710 1.280 ;
        RECT 885.830 0.270 890.230 1.280 ;
        RECT 891.350 0.270 895.750 1.280 ;
        RECT 896.870 0.270 901.270 1.280 ;
        RECT 902.390 0.270 906.790 1.280 ;
        RECT 907.910 0.270 912.310 1.280 ;
        RECT 913.430 0.270 917.830 1.280 ;
        RECT 918.950 0.270 923.350 1.280 ;
        RECT 924.470 0.270 928.870 1.280 ;
        RECT 929.990 0.270 934.390 1.280 ;
        RECT 935.510 0.270 939.910 1.280 ;
        RECT 941.030 0.270 945.430 1.280 ;
        RECT 946.550 0.270 950.950 1.280 ;
        RECT 952.070 0.270 956.470 1.280 ;
        RECT 957.590 0.270 961.990 1.280 ;
        RECT 963.110 0.270 967.510 1.280 ;
        RECT 968.630 0.270 973.030 1.280 ;
        RECT 974.150 0.270 978.550 1.280 ;
        RECT 979.670 0.270 984.070 1.280 ;
        RECT 985.190 0.270 989.590 1.280 ;
        RECT 990.710 0.270 995.110 1.280 ;
        RECT 996.230 0.270 1000.630 1.280 ;
        RECT 1001.750 0.270 1006.150 1.280 ;
        RECT 1007.270 0.270 1011.670 1.280 ;
        RECT 1012.790 0.270 1017.190 1.280 ;
        RECT 1018.310 0.270 1022.710 1.280 ;
        RECT 1023.830 0.270 1028.230 1.280 ;
        RECT 1029.350 0.270 1033.750 1.280 ;
        RECT 1034.870 0.270 1039.270 1.280 ;
        RECT 1040.390 0.270 1044.790 1.280 ;
        RECT 1045.910 0.270 1050.310 1.280 ;
        RECT 1051.430 0.270 1055.830 1.280 ;
        RECT 1056.950 0.270 1061.350 1.280 ;
        RECT 1062.470 0.270 1066.870 1.280 ;
        RECT 1067.990 0.270 1072.390 1.280 ;
        RECT 1073.510 0.270 1077.910 1.280 ;
        RECT 1079.030 0.270 1083.430 1.280 ;
        RECT 1084.550 0.270 1088.950 1.280 ;
        RECT 1090.070 0.270 1094.470 1.280 ;
        RECT 1095.590 0.270 1099.990 1.280 ;
        RECT 1101.110 0.270 1105.510 1.280 ;
        RECT 1106.630 0.270 1111.030 1.280 ;
        RECT 1112.150 0.270 1116.550 1.280 ;
        RECT 1117.670 0.270 1122.070 1.280 ;
        RECT 1123.190 0.270 1127.590 1.280 ;
        RECT 1128.710 0.270 1133.110 1.280 ;
        RECT 1134.230 0.270 1138.630 1.280 ;
        RECT 1139.750 0.270 1144.150 1.280 ;
        RECT 1145.270 0.270 1149.670 1.280 ;
        RECT 1150.790 0.270 1155.190 1.280 ;
        RECT 1156.310 0.270 1160.710 1.280 ;
        RECT 1161.830 0.270 1166.230 1.280 ;
        RECT 1167.350 0.270 1171.750 1.280 ;
        RECT 1172.870 0.270 1177.270 1.280 ;
        RECT 1178.390 0.270 1182.790 1.280 ;
        RECT 1183.910 0.270 1188.310 1.280 ;
        RECT 1189.430 0.270 1193.830 1.280 ;
        RECT 1194.950 0.270 1199.350 1.280 ;
        RECT 1200.470 0.270 1204.870 1.280 ;
        RECT 1205.990 0.270 1210.390 1.280 ;
        RECT 1211.510 0.270 1215.910 1.280 ;
        RECT 1217.030 0.270 1221.430 1.280 ;
        RECT 1222.550 0.270 1226.950 1.280 ;
        RECT 1228.070 0.270 1232.470 1.280 ;
        RECT 1233.590 0.270 1237.990 1.280 ;
        RECT 1239.110 0.270 1243.510 1.280 ;
        RECT 1244.630 0.270 1249.030 1.280 ;
        RECT 1250.150 0.270 1254.550 1.280 ;
        RECT 1255.670 0.270 1260.070 1.280 ;
        RECT 1261.190 0.270 1265.590 1.280 ;
        RECT 1266.710 0.270 1271.110 1.280 ;
        RECT 1272.230 0.270 1276.630 1.280 ;
        RECT 1277.750 0.270 1282.150 1.280 ;
        RECT 1283.270 0.270 1287.670 1.280 ;
        RECT 1288.790 0.270 1293.190 1.280 ;
        RECT 1294.310 0.270 1298.710 1.280 ;
        RECT 1299.830 0.270 1304.230 1.280 ;
        RECT 1305.350 0.270 1309.750 1.280 ;
        RECT 1310.870 0.270 1315.270 1.280 ;
        RECT 1316.390 0.270 1320.790 1.280 ;
        RECT 1321.910 0.270 1326.310 1.280 ;
        RECT 1327.430 0.270 1331.830 1.280 ;
        RECT 1332.950 0.270 1337.350 1.280 ;
        RECT 1338.470 0.270 1342.870 1.280 ;
        RECT 1343.990 0.270 1348.390 1.280 ;
        RECT 1349.510 0.270 1353.910 1.280 ;
        RECT 1355.030 0.270 1359.430 1.280 ;
        RECT 1360.550 0.270 1364.950 1.280 ;
        RECT 1366.070 0.270 1370.470 1.280 ;
        RECT 1371.590 0.270 1375.990 1.280 ;
        RECT 1377.110 0.270 1381.510 1.280 ;
        RECT 1382.630 0.270 1387.030 1.280 ;
        RECT 1388.150 0.270 1392.550 1.280 ;
        RECT 1393.670 0.270 1398.070 1.280 ;
        RECT 1399.190 0.270 1403.590 1.280 ;
        RECT 1404.710 0.270 1409.110 1.280 ;
        RECT 1410.230 0.270 1414.630 1.280 ;
        RECT 1415.750 0.270 1420.150 1.280 ;
        RECT 1421.270 0.270 1425.670 1.280 ;
        RECT 1426.790 0.270 1431.190 1.280 ;
        RECT 1432.310 0.270 1436.710 1.280 ;
        RECT 1437.830 0.270 1442.230 1.280 ;
        RECT 1443.350 0.270 1447.750 1.280 ;
        RECT 1448.870 0.270 1453.270 1.280 ;
        RECT 1454.390 0.270 1458.790 1.280 ;
        RECT 1459.910 0.270 1464.310 1.280 ;
        RECT 1465.430 0.270 1469.830 1.280 ;
        RECT 1470.950 0.270 1475.350 1.280 ;
        RECT 1476.470 0.270 1480.870 1.280 ;
        RECT 1481.990 0.270 1486.390 1.280 ;
        RECT 1487.510 0.270 1491.910 1.280 ;
        RECT 1493.030 0.270 1497.430 1.280 ;
        RECT 1498.550 0.270 1502.950 1.280 ;
        RECT 1504.070 0.270 1508.470 1.280 ;
        RECT 1509.590 0.270 1513.990 1.280 ;
        RECT 1515.110 0.270 1519.510 1.280 ;
        RECT 1520.630 0.270 1525.030 1.280 ;
        RECT 1526.150 0.270 1530.550 1.280 ;
        RECT 1531.670 0.270 1536.070 1.280 ;
        RECT 1537.190 0.270 1541.590 1.280 ;
        RECT 1542.710 0.270 1547.110 1.280 ;
        RECT 1548.230 0.270 1552.630 1.280 ;
        RECT 1553.750 0.270 1558.150 1.280 ;
        RECT 1559.270 0.270 1563.670 1.280 ;
        RECT 1564.790 0.270 1569.190 1.280 ;
        RECT 1570.310 0.270 1574.710 1.280 ;
        RECT 1575.830 0.270 1580.230 1.280 ;
        RECT 1581.350 0.270 1585.750 1.280 ;
        RECT 1586.870 0.270 1591.270 1.280 ;
        RECT 1592.390 0.270 1596.790 1.280 ;
        RECT 1597.910 0.270 1602.310 1.280 ;
        RECT 1603.430 0.270 1607.830 1.280 ;
        RECT 1608.950 0.270 1613.350 1.280 ;
        RECT 1614.470 0.270 1618.870 1.280 ;
        RECT 1619.990 0.270 1624.390 1.280 ;
        RECT 1625.510 0.270 1629.910 1.280 ;
        RECT 1631.030 0.270 1635.430 1.280 ;
        RECT 1636.550 0.270 1640.950 1.280 ;
        RECT 1642.070 0.270 1646.470 1.280 ;
        RECT 1647.590 0.270 1651.990 1.280 ;
        RECT 1653.110 0.270 1657.510 1.280 ;
        RECT 1658.630 0.270 1663.030 1.280 ;
        RECT 1664.150 0.270 1668.550 1.280 ;
        RECT 1669.670 0.270 1674.070 1.280 ;
        RECT 1675.190 0.270 1679.590 1.280 ;
        RECT 1680.710 0.270 1685.110 1.280 ;
        RECT 1686.230 0.270 1690.630 1.280 ;
        RECT 1691.750 0.270 1696.150 1.280 ;
        RECT 1697.270 0.270 1701.670 1.280 ;
        RECT 1702.790 0.270 1707.190 1.280 ;
        RECT 1708.310 0.270 1712.710 1.280 ;
        RECT 1713.830 0.270 1718.230 1.280 ;
        RECT 1719.350 0.270 1723.750 1.280 ;
        RECT 1724.870 0.270 1729.270 1.280 ;
        RECT 1730.390 0.270 1734.790 1.280 ;
        RECT 1735.910 0.270 1740.310 1.280 ;
        RECT 1741.430 0.270 1745.830 1.280 ;
        RECT 1746.950 0.270 1751.350 1.280 ;
        RECT 1752.470 0.270 1756.870 1.280 ;
        RECT 1757.990 0.270 1762.390 1.280 ;
        RECT 1763.510 0.270 1767.910 1.280 ;
        RECT 1769.030 0.270 1773.430 1.280 ;
        RECT 1774.550 0.270 1778.950 1.280 ;
        RECT 1780.070 0.270 1784.470 1.280 ;
        RECT 1785.590 0.270 1789.990 1.280 ;
        RECT 1791.110 0.270 1795.510 1.280 ;
        RECT 1796.630 0.270 1801.030 1.280 ;
        RECT 1802.150 0.270 1806.550 1.280 ;
        RECT 1807.670 0.270 1812.070 1.280 ;
        RECT 1813.190 0.270 1817.590 1.280 ;
        RECT 1818.710 0.270 1823.110 1.280 ;
        RECT 1824.230 0.270 1828.630 1.280 ;
        RECT 1829.750 0.270 1834.150 1.280 ;
        RECT 1835.270 0.270 1839.670 1.280 ;
        RECT 1840.790 0.270 1845.190 1.280 ;
        RECT 1846.310 0.270 1850.710 1.280 ;
        RECT 1851.830 0.270 1856.230 1.280 ;
        RECT 1857.350 0.270 1861.750 1.280 ;
        RECT 1862.870 0.270 1867.270 1.280 ;
        RECT 1868.390 0.270 1872.790 1.280 ;
        RECT 1873.910 0.270 1878.310 1.280 ;
        RECT 1879.430 0.270 1883.830 1.280 ;
        RECT 1884.950 0.270 1889.350 1.280 ;
        RECT 1890.470 0.270 1894.870 1.280 ;
        RECT 1895.990 0.270 1900.390 1.280 ;
        RECT 1901.510 0.270 1905.910 1.280 ;
        RECT 1907.030 0.270 1911.430 1.280 ;
        RECT 1912.550 0.270 1916.950 1.280 ;
        RECT 1918.070 0.270 1922.470 1.280 ;
        RECT 1923.590 0.270 1927.990 1.280 ;
        RECT 1929.110 0.270 1933.510 1.280 ;
        RECT 1934.630 0.270 1939.030 1.280 ;
        RECT 1940.150 0.270 1944.550 1.280 ;
        RECT 1945.670 0.270 1950.070 1.280 ;
        RECT 1951.190 0.270 1955.590 1.280 ;
        RECT 1956.710 0.270 1961.110 1.280 ;
        RECT 1962.230 0.270 1966.630 1.280 ;
        RECT 1967.750 0.270 1972.150 1.280 ;
        RECT 1973.270 0.270 1977.670 1.280 ;
        RECT 1978.790 0.270 1983.190 1.280 ;
        RECT 1984.310 0.270 1988.710 1.280 ;
        RECT 1989.830 0.270 1994.230 1.280 ;
        RECT 1995.350 0.270 1999.750 1.280 ;
        RECT 2000.870 0.270 2005.270 1.280 ;
        RECT 2006.390 0.270 2010.790 1.280 ;
        RECT 2011.910 0.270 2016.310 1.280 ;
        RECT 2017.430 0.270 2021.830 1.280 ;
        RECT 2022.950 0.270 2027.350 1.280 ;
        RECT 2028.470 0.270 2032.870 1.280 ;
        RECT 2033.990 0.270 2038.390 1.280 ;
        RECT 2039.510 0.270 2043.910 1.280 ;
        RECT 2045.030 0.270 2049.430 1.280 ;
        RECT 2050.550 0.270 2054.950 1.280 ;
        RECT 2056.070 0.270 2060.470 1.280 ;
        RECT 2061.590 0.270 2065.990 1.280 ;
        RECT 2067.110 0.270 2071.510 1.280 ;
        RECT 2072.630 0.270 2077.030 1.280 ;
        RECT 2078.150 0.270 2082.550 1.280 ;
        RECT 2083.670 0.270 2088.070 1.280 ;
        RECT 2089.190 0.270 2093.590 1.280 ;
        RECT 2094.710 0.270 2099.110 1.280 ;
        RECT 2100.230 0.270 2104.630 1.280 ;
        RECT 2105.750 0.270 2110.150 1.280 ;
        RECT 2111.270 0.270 2115.670 1.280 ;
        RECT 2116.790 0.270 2121.190 1.280 ;
        RECT 2122.310 0.270 2126.710 1.280 ;
        RECT 2127.830 0.270 2132.230 1.280 ;
        RECT 2133.350 0.270 2137.750 1.280 ;
        RECT 2138.870 0.270 2143.270 1.280 ;
        RECT 2144.390 0.270 2148.790 1.280 ;
        RECT 2149.910 0.270 2154.310 1.280 ;
        RECT 2155.430 0.270 2159.830 1.280 ;
        RECT 2160.950 0.270 2165.350 1.280 ;
        RECT 2166.470 0.270 2170.870 1.280 ;
        RECT 2171.990 0.270 2176.390 1.280 ;
        RECT 2177.510 0.270 2181.910 1.280 ;
        RECT 2183.030 0.270 2187.430 1.280 ;
        RECT 2188.550 0.270 2192.950 1.280 ;
        RECT 2194.070 0.270 2198.470 1.280 ;
        RECT 2199.590 0.270 2203.990 1.280 ;
        RECT 2205.110 0.270 2209.510 1.280 ;
        RECT 2210.630 0.270 2215.030 1.280 ;
        RECT 2216.150 0.270 2220.550 1.280 ;
        RECT 2221.670 0.270 2226.070 1.280 ;
        RECT 2227.190 0.270 2231.590 1.280 ;
        RECT 2232.710 0.270 2237.110 1.280 ;
        RECT 2238.230 0.270 2242.630 1.280 ;
        RECT 2243.750 0.270 2248.150 1.280 ;
        RECT 2249.270 0.270 2253.670 1.280 ;
        RECT 2254.790 0.270 2259.190 1.280 ;
        RECT 2260.310 0.270 2264.710 1.280 ;
        RECT 2265.830 0.270 2270.230 1.280 ;
        RECT 2271.350 0.270 2275.750 1.280 ;
        RECT 2276.870 0.270 2281.270 1.280 ;
        RECT 2282.390 0.270 2286.790 1.280 ;
        RECT 2287.910 0.270 2292.310 1.280 ;
        RECT 2293.430 0.270 2297.830 1.280 ;
        RECT 2298.950 0.270 2303.350 1.280 ;
        RECT 2304.470 0.270 2308.870 1.280 ;
        RECT 2309.990 0.270 2314.390 1.280 ;
        RECT 2315.510 0.270 2319.910 1.280 ;
        RECT 2321.030 0.270 2325.430 1.280 ;
        RECT 2326.550 0.270 2330.950 1.280 ;
        RECT 2332.070 0.270 2336.470 1.280 ;
        RECT 2337.590 0.270 2341.990 1.280 ;
        RECT 2343.110 0.270 2347.510 1.280 ;
        RECT 2348.630 0.270 2353.030 1.280 ;
        RECT 2354.150 0.270 2358.550 1.280 ;
        RECT 2359.670 0.270 2364.070 1.280 ;
        RECT 2365.190 0.270 2369.590 1.280 ;
        RECT 2370.710 0.270 2375.110 1.280 ;
        RECT 2376.230 0.270 2380.630 1.280 ;
        RECT 2381.750 0.270 2386.150 1.280 ;
        RECT 2387.270 0.270 2391.670 1.280 ;
        RECT 2392.790 0.270 2397.190 1.280 ;
        RECT 2398.310 0.270 2402.710 1.280 ;
        RECT 2403.830 0.270 2408.230 1.280 ;
        RECT 2409.350 0.270 2413.750 1.280 ;
        RECT 2414.870 0.270 2419.270 1.280 ;
        RECT 2420.390 0.270 2424.790 1.280 ;
        RECT 2425.910 0.270 2430.310 1.280 ;
        RECT 2431.430 0.270 2435.830 1.280 ;
        RECT 2436.950 0.270 2441.350 1.280 ;
        RECT 2442.470 0.270 2446.870 1.280 ;
        RECT 2447.990 0.270 2452.390 1.280 ;
        RECT 2453.510 0.270 2457.910 1.280 ;
        RECT 2459.030 0.270 2463.430 1.280 ;
        RECT 2464.550 0.270 2468.950 1.280 ;
        RECT 2470.070 0.270 2474.470 1.280 ;
        RECT 2475.590 0.270 2479.990 1.280 ;
        RECT 2481.110 0.270 2485.510 1.280 ;
        RECT 2486.630 0.270 2491.030 1.280 ;
        RECT 2492.150 0.270 2496.550 1.280 ;
        RECT 2497.670 0.270 2502.070 1.280 ;
        RECT 2503.190 0.270 2507.590 1.280 ;
        RECT 2508.710 0.270 2513.110 1.280 ;
        RECT 2514.230 0.270 2518.630 1.280 ;
        RECT 2519.750 0.270 2524.150 1.280 ;
        RECT 2525.270 0.270 2529.670 1.280 ;
        RECT 2530.790 0.270 2535.190 1.280 ;
        RECT 2536.310 0.270 2540.710 1.280 ;
        RECT 2541.830 0.270 2546.230 1.280 ;
        RECT 2547.350 0.270 2551.750 1.280 ;
        RECT 2552.870 0.270 2557.270 1.280 ;
        RECT 2558.390 0.270 2562.790 1.280 ;
        RECT 2563.910 0.270 2568.310 1.280 ;
        RECT 2569.430 0.270 2573.830 1.280 ;
        RECT 2574.950 0.270 2579.350 1.280 ;
        RECT 2580.470 0.270 2584.870 1.280 ;
        RECT 2585.990 0.270 2590.390 1.280 ;
        RECT 2591.510 0.270 2595.910 1.280 ;
        RECT 2597.030 0.270 2601.430 1.280 ;
        RECT 2602.550 0.270 2606.950 1.280 ;
        RECT 2608.070 0.270 2612.470 1.280 ;
        RECT 2613.590 0.270 2617.990 1.280 ;
        RECT 2619.110 0.270 2623.510 1.280 ;
        RECT 2624.630 0.270 2629.030 1.280 ;
        RECT 2630.150 0.270 2634.550 1.280 ;
        RECT 2635.670 0.270 2640.070 1.280 ;
        RECT 2641.190 0.270 2645.590 1.280 ;
        RECT 2646.710 0.270 2651.110 1.280 ;
        RECT 2652.230 0.270 2656.630 1.280 ;
        RECT 2657.750 0.270 2662.150 1.280 ;
        RECT 2663.270 0.270 2667.670 1.280 ;
        RECT 2668.790 0.270 2673.190 1.280 ;
        RECT 2674.310 0.270 2678.710 1.280 ;
        RECT 2679.830 0.270 2684.230 1.280 ;
        RECT 2685.350 0.270 2689.750 1.280 ;
        RECT 2690.870 0.270 2695.270 1.280 ;
        RECT 2696.390 0.270 2700.790 1.280 ;
        RECT 2701.910 0.270 2706.310 1.280 ;
        RECT 2707.430 0.270 2711.830 1.280 ;
        RECT 2712.950 0.270 2717.350 1.280 ;
        RECT 2718.470 0.270 2722.870 1.280 ;
        RECT 2723.990 0.270 2728.390 1.280 ;
        RECT 2729.510 0.270 2733.910 1.280 ;
        RECT 2735.030 0.270 2739.430 1.280 ;
        RECT 2740.550 0.270 2744.950 1.280 ;
        RECT 2746.070 0.270 2750.470 1.280 ;
        RECT 2751.590 0.270 2755.990 1.280 ;
        RECT 2757.110 0.270 2761.510 1.280 ;
        RECT 2762.630 0.270 2767.030 1.280 ;
        RECT 2768.150 0.270 2772.550 1.280 ;
        RECT 2773.670 0.270 2778.070 1.280 ;
        RECT 2779.190 0.270 2783.590 1.280 ;
        RECT 2784.710 0.270 2789.110 1.280 ;
        RECT 2790.230 0.270 2794.630 1.280 ;
        RECT 2795.750 0.270 2800.150 1.280 ;
        RECT 2801.270 0.270 2871.690 1.280 ;
      LAYER met3 ;
        RECT 1.000 3438.060 2879.000 3468.165 ;
        RECT 1.000 3436.060 2878.600 3438.060 ;
        RECT 1.000 3434.660 2879.000 3436.060 ;
        RECT 1.400 3432.660 2879.000 3434.660 ;
        RECT 1.000 3372.780 2879.000 3432.660 ;
        RECT 1.000 3370.780 2878.600 3372.780 ;
        RECT 1.000 3370.740 2879.000 3370.780 ;
        RECT 1.400 3368.740 2879.000 3370.740 ;
        RECT 1.000 3307.500 2879.000 3368.740 ;
        RECT 1.000 3306.820 2878.600 3307.500 ;
        RECT 1.400 3305.500 2878.600 3306.820 ;
        RECT 1.400 3304.820 2879.000 3305.500 ;
        RECT 1.000 3242.900 2879.000 3304.820 ;
        RECT 1.400 3242.220 2879.000 3242.900 ;
        RECT 1.400 3240.900 2878.600 3242.220 ;
        RECT 1.000 3240.220 2878.600 3240.900 ;
        RECT 1.000 3178.980 2879.000 3240.220 ;
        RECT 1.400 3176.980 2879.000 3178.980 ;
        RECT 1.000 3176.940 2879.000 3176.980 ;
        RECT 1.000 3174.940 2878.600 3176.940 ;
        RECT 1.000 3115.060 2879.000 3174.940 ;
        RECT 1.400 3113.060 2879.000 3115.060 ;
        RECT 1.000 3111.660 2879.000 3113.060 ;
        RECT 1.000 3109.660 2878.600 3111.660 ;
        RECT 1.000 3051.140 2879.000 3109.660 ;
        RECT 1.400 3049.140 2879.000 3051.140 ;
        RECT 1.000 3046.380 2879.000 3049.140 ;
        RECT 1.000 3044.380 2878.600 3046.380 ;
        RECT 1.000 2987.220 2879.000 3044.380 ;
        RECT 1.400 2985.220 2879.000 2987.220 ;
        RECT 1.000 2981.100 2879.000 2985.220 ;
        RECT 1.000 2979.100 2878.600 2981.100 ;
        RECT 1.000 2923.300 2879.000 2979.100 ;
        RECT 1.400 2921.300 2879.000 2923.300 ;
        RECT 1.000 2915.820 2879.000 2921.300 ;
        RECT 1.000 2913.820 2878.600 2915.820 ;
        RECT 1.000 2859.380 2879.000 2913.820 ;
        RECT 1.400 2857.380 2879.000 2859.380 ;
        RECT 1.000 2850.540 2879.000 2857.380 ;
        RECT 1.000 2848.540 2878.600 2850.540 ;
        RECT 1.000 2795.460 2879.000 2848.540 ;
        RECT 1.400 2793.460 2879.000 2795.460 ;
        RECT 1.000 2785.260 2879.000 2793.460 ;
        RECT 1.000 2783.260 2878.600 2785.260 ;
        RECT 1.000 2731.540 2879.000 2783.260 ;
        RECT 1.400 2729.540 2879.000 2731.540 ;
        RECT 1.000 2719.980 2879.000 2729.540 ;
        RECT 1.000 2717.980 2878.600 2719.980 ;
        RECT 1.000 2667.620 2879.000 2717.980 ;
        RECT 1.400 2665.620 2879.000 2667.620 ;
        RECT 1.000 2654.700 2879.000 2665.620 ;
        RECT 1.000 2652.700 2878.600 2654.700 ;
        RECT 1.000 2603.700 2879.000 2652.700 ;
        RECT 1.400 2601.700 2879.000 2603.700 ;
        RECT 1.000 2589.420 2879.000 2601.700 ;
        RECT 1.000 2587.420 2878.600 2589.420 ;
        RECT 1.000 2539.780 2879.000 2587.420 ;
        RECT 1.400 2537.780 2879.000 2539.780 ;
        RECT 1.000 2524.140 2879.000 2537.780 ;
        RECT 1.000 2522.140 2878.600 2524.140 ;
        RECT 1.000 2475.860 2879.000 2522.140 ;
        RECT 1.400 2473.860 2879.000 2475.860 ;
        RECT 1.000 2458.860 2879.000 2473.860 ;
        RECT 1.000 2456.860 2878.600 2458.860 ;
        RECT 1.000 2411.940 2879.000 2456.860 ;
        RECT 1.400 2409.940 2879.000 2411.940 ;
        RECT 1.000 2393.580 2879.000 2409.940 ;
        RECT 1.000 2391.580 2878.600 2393.580 ;
        RECT 1.000 2348.020 2879.000 2391.580 ;
        RECT 1.400 2346.020 2879.000 2348.020 ;
        RECT 1.000 2328.300 2879.000 2346.020 ;
        RECT 1.000 2326.300 2878.600 2328.300 ;
        RECT 1.000 2284.100 2879.000 2326.300 ;
        RECT 1.400 2282.100 2879.000 2284.100 ;
        RECT 1.000 2263.020 2879.000 2282.100 ;
        RECT 1.000 2261.020 2878.600 2263.020 ;
        RECT 1.000 2220.180 2879.000 2261.020 ;
        RECT 1.400 2218.180 2879.000 2220.180 ;
        RECT 1.000 2197.740 2879.000 2218.180 ;
        RECT 1.000 2195.740 2878.600 2197.740 ;
        RECT 1.000 2156.260 2879.000 2195.740 ;
        RECT 1.400 2154.260 2879.000 2156.260 ;
        RECT 1.000 2132.460 2879.000 2154.260 ;
        RECT 1.000 2130.460 2878.600 2132.460 ;
        RECT 1.000 2092.340 2879.000 2130.460 ;
        RECT 1.400 2090.340 2879.000 2092.340 ;
        RECT 1.000 2067.180 2879.000 2090.340 ;
        RECT 1.000 2065.180 2878.600 2067.180 ;
        RECT 1.000 2028.420 2879.000 2065.180 ;
        RECT 1.400 2026.420 2879.000 2028.420 ;
        RECT 1.000 2001.900 2879.000 2026.420 ;
        RECT 1.000 1999.900 2878.600 2001.900 ;
        RECT 1.000 1964.500 2879.000 1999.900 ;
        RECT 1.400 1962.500 2879.000 1964.500 ;
        RECT 1.000 1936.620 2879.000 1962.500 ;
        RECT 1.000 1934.620 2878.600 1936.620 ;
        RECT 1.000 1900.580 2879.000 1934.620 ;
        RECT 1.400 1898.580 2879.000 1900.580 ;
        RECT 1.000 1871.340 2879.000 1898.580 ;
        RECT 1.000 1869.340 2878.600 1871.340 ;
        RECT 1.000 1836.660 2879.000 1869.340 ;
        RECT 1.400 1834.660 2879.000 1836.660 ;
        RECT 1.000 1806.060 2879.000 1834.660 ;
        RECT 1.000 1804.060 2878.600 1806.060 ;
        RECT 1.000 1772.740 2879.000 1804.060 ;
        RECT 1.400 1770.740 2879.000 1772.740 ;
        RECT 1.000 1740.780 2879.000 1770.740 ;
        RECT 1.000 1738.780 2878.600 1740.780 ;
        RECT 1.000 1708.820 2879.000 1738.780 ;
        RECT 1.400 1706.820 2879.000 1708.820 ;
        RECT 1.000 1675.500 2879.000 1706.820 ;
        RECT 1.000 1673.500 2878.600 1675.500 ;
        RECT 1.000 1644.900 2879.000 1673.500 ;
        RECT 1.400 1642.900 2879.000 1644.900 ;
        RECT 1.000 1610.220 2879.000 1642.900 ;
        RECT 1.000 1608.220 2878.600 1610.220 ;
        RECT 1.000 1580.980 2879.000 1608.220 ;
        RECT 1.400 1578.980 2879.000 1580.980 ;
        RECT 1.000 1544.940 2879.000 1578.980 ;
        RECT 1.000 1542.940 2878.600 1544.940 ;
        RECT 1.000 1517.060 2879.000 1542.940 ;
        RECT 1.400 1515.060 2879.000 1517.060 ;
        RECT 1.000 1479.660 2879.000 1515.060 ;
        RECT 1.000 1477.660 2878.600 1479.660 ;
        RECT 1.000 1453.140 2879.000 1477.660 ;
        RECT 1.400 1451.140 2879.000 1453.140 ;
        RECT 1.000 1414.380 2879.000 1451.140 ;
        RECT 1.000 1412.380 2878.600 1414.380 ;
        RECT 1.000 1389.220 2879.000 1412.380 ;
        RECT 1.400 1387.220 2879.000 1389.220 ;
        RECT 1.000 1349.100 2879.000 1387.220 ;
        RECT 1.000 1347.100 2878.600 1349.100 ;
        RECT 1.000 1325.300 2879.000 1347.100 ;
        RECT 1.400 1323.300 2879.000 1325.300 ;
        RECT 1.000 1283.820 2879.000 1323.300 ;
        RECT 1.000 1281.820 2878.600 1283.820 ;
        RECT 1.000 1261.380 2879.000 1281.820 ;
        RECT 1.400 1259.380 2879.000 1261.380 ;
        RECT 1.000 1218.540 2879.000 1259.380 ;
        RECT 1.000 1216.540 2878.600 1218.540 ;
        RECT 1.000 1197.460 2879.000 1216.540 ;
        RECT 1.400 1195.460 2879.000 1197.460 ;
        RECT 1.000 1153.260 2879.000 1195.460 ;
        RECT 1.000 1151.260 2878.600 1153.260 ;
        RECT 1.000 1133.540 2879.000 1151.260 ;
        RECT 1.400 1131.540 2879.000 1133.540 ;
        RECT 1.000 1087.980 2879.000 1131.540 ;
        RECT 1.000 1085.980 2878.600 1087.980 ;
        RECT 1.000 1069.620 2879.000 1085.980 ;
        RECT 1.400 1067.620 2879.000 1069.620 ;
        RECT 1.000 1022.700 2879.000 1067.620 ;
        RECT 1.000 1020.700 2878.600 1022.700 ;
        RECT 1.000 1005.700 2879.000 1020.700 ;
        RECT 1.400 1003.700 2879.000 1005.700 ;
        RECT 1.000 957.420 2879.000 1003.700 ;
        RECT 1.000 955.420 2878.600 957.420 ;
        RECT 1.000 941.780 2879.000 955.420 ;
        RECT 1.400 939.780 2879.000 941.780 ;
        RECT 1.000 892.140 2879.000 939.780 ;
        RECT 1.000 890.140 2878.600 892.140 ;
        RECT 1.000 877.860 2879.000 890.140 ;
        RECT 1.400 875.860 2879.000 877.860 ;
        RECT 1.000 826.860 2879.000 875.860 ;
        RECT 1.000 824.860 2878.600 826.860 ;
        RECT 1.000 813.940 2879.000 824.860 ;
        RECT 1.400 811.940 2879.000 813.940 ;
        RECT 1.000 761.580 2879.000 811.940 ;
        RECT 1.000 759.580 2878.600 761.580 ;
        RECT 1.000 750.020 2879.000 759.580 ;
        RECT 1.400 748.020 2879.000 750.020 ;
        RECT 1.000 696.300 2879.000 748.020 ;
        RECT 1.000 694.300 2878.600 696.300 ;
        RECT 1.000 686.100 2879.000 694.300 ;
        RECT 1.400 684.100 2879.000 686.100 ;
        RECT 1.000 631.020 2879.000 684.100 ;
        RECT 1.000 629.020 2878.600 631.020 ;
        RECT 1.000 622.180 2879.000 629.020 ;
        RECT 1.400 620.180 2879.000 622.180 ;
        RECT 1.000 565.740 2879.000 620.180 ;
        RECT 1.000 563.740 2878.600 565.740 ;
        RECT 1.000 558.260 2879.000 563.740 ;
        RECT 1.400 556.260 2879.000 558.260 ;
        RECT 1.000 500.460 2879.000 556.260 ;
        RECT 1.000 498.460 2878.600 500.460 ;
        RECT 1.000 494.340 2879.000 498.460 ;
        RECT 1.400 492.340 2879.000 494.340 ;
        RECT 1.000 435.180 2879.000 492.340 ;
        RECT 1.000 433.180 2878.600 435.180 ;
        RECT 1.000 430.420 2879.000 433.180 ;
        RECT 1.400 428.420 2879.000 430.420 ;
        RECT 1.000 369.900 2879.000 428.420 ;
        RECT 1.000 367.900 2878.600 369.900 ;
        RECT 1.000 366.500 2879.000 367.900 ;
        RECT 1.400 364.500 2879.000 366.500 ;
        RECT 1.000 304.620 2879.000 364.500 ;
        RECT 1.000 302.620 2878.600 304.620 ;
        RECT 1.000 302.580 2879.000 302.620 ;
        RECT 1.400 300.580 2879.000 302.580 ;
        RECT 1.000 239.340 2879.000 300.580 ;
        RECT 1.000 238.660 2878.600 239.340 ;
        RECT 1.400 237.340 2878.600 238.660 ;
        RECT 1.400 236.660 2879.000 237.340 ;
        RECT 1.000 174.740 2879.000 236.660 ;
        RECT 1.400 174.060 2879.000 174.740 ;
        RECT 1.400 172.740 2878.600 174.060 ;
        RECT 1.000 172.060 2878.600 172.740 ;
        RECT 1.000 110.820 2879.000 172.060 ;
        RECT 1.400 108.820 2879.000 110.820 ;
        RECT 1.000 108.780 2879.000 108.820 ;
        RECT 1.000 106.780 2878.600 108.780 ;
        RECT 1.000 46.900 2879.000 106.780 ;
        RECT 1.400 44.900 2879.000 46.900 ;
        RECT 1.000 43.500 2879.000 44.900 ;
        RECT 1.000 41.500 2878.600 43.500 ;
        RECT 1.000 6.975 2879.000 41.500 ;
      LAYER met4 ;
        RECT 53.655 3411.140 98.570 3467.145 ;
        RECT 102.470 3411.140 188.570 3467.145 ;
        RECT 192.470 3411.140 278.570 3467.145 ;
        RECT 282.470 3411.140 368.570 3467.145 ;
        RECT 372.470 3411.140 458.570 3467.145 ;
        RECT 462.470 3411.140 548.570 3467.145 ;
        RECT 552.470 3411.140 638.570 3467.145 ;
        RECT 642.470 3411.140 728.570 3467.145 ;
        RECT 732.470 3411.140 818.570 3467.145 ;
        RECT 53.655 2975.400 818.570 3411.140 ;
        RECT 53.655 2851.140 98.570 2975.400 ;
        RECT 102.470 2851.140 188.570 2975.400 ;
        RECT 192.470 2851.140 278.570 2975.400 ;
        RECT 282.470 2851.140 368.570 2975.400 ;
        RECT 372.470 2851.140 458.570 2975.400 ;
        RECT 462.470 2851.140 548.570 2975.400 ;
        RECT 552.470 2851.140 638.570 2975.400 ;
        RECT 642.470 2851.140 728.570 2975.400 ;
        RECT 732.470 2851.140 818.570 2975.400 ;
        RECT 53.655 2415.400 818.570 2851.140 ;
        RECT 53.655 2256.140 98.570 2415.400 ;
        RECT 102.470 2256.140 188.570 2415.400 ;
        RECT 192.470 2256.140 278.570 2415.400 ;
        RECT 282.470 2256.140 368.570 2415.400 ;
        RECT 372.470 2256.140 458.570 2415.400 ;
        RECT 462.470 2256.140 548.570 2415.400 ;
        RECT 552.470 2256.140 638.570 2415.400 ;
        RECT 642.470 2256.140 728.570 2415.400 ;
        RECT 732.470 2256.140 818.570 2415.400 ;
        RECT 53.655 1820.400 818.570 2256.140 ;
        RECT 53.655 1696.140 98.570 1820.400 ;
        RECT 102.470 1696.140 188.570 1820.400 ;
        RECT 192.470 1696.140 278.570 1820.400 ;
        RECT 282.470 1696.140 368.570 1820.400 ;
        RECT 372.470 1696.140 458.570 1820.400 ;
        RECT 462.470 1696.140 548.570 1820.400 ;
        RECT 552.470 1696.140 638.570 1820.400 ;
        RECT 642.470 1696.140 728.570 1820.400 ;
        RECT 732.470 1696.140 818.570 1820.400 ;
        RECT 53.655 1260.400 818.570 1696.140 ;
        RECT 53.655 1116.140 98.570 1260.400 ;
        RECT 102.470 1116.140 188.570 1260.400 ;
        RECT 192.470 1116.140 278.570 1260.400 ;
        RECT 282.470 1116.140 368.570 1260.400 ;
        RECT 372.470 1116.140 458.570 1260.400 ;
        RECT 462.470 1116.140 548.570 1260.400 ;
        RECT 552.470 1116.140 638.570 1260.400 ;
        RECT 642.470 1116.140 728.570 1260.400 ;
        RECT 732.470 1116.140 818.570 1260.400 ;
        RECT 53.655 680.400 818.570 1116.140 ;
        RECT 53.655 551.140 98.570 680.400 ;
        RECT 102.470 551.140 188.570 680.400 ;
        RECT 192.470 551.140 278.570 680.400 ;
        RECT 282.470 551.140 368.570 680.400 ;
        RECT 372.470 551.140 458.570 680.400 ;
        RECT 462.470 551.140 548.570 680.400 ;
        RECT 552.470 551.140 638.570 680.400 ;
        RECT 642.470 551.140 728.570 680.400 ;
        RECT 732.470 551.140 818.570 680.400 ;
        RECT 53.655 115.400 818.570 551.140 ;
        RECT 53.655 10.240 98.570 115.400 ;
        RECT 102.470 10.240 188.570 115.400 ;
        RECT 192.470 10.240 278.570 115.400 ;
        RECT 282.470 10.240 368.570 115.400 ;
        RECT 372.470 10.240 458.570 115.400 ;
        RECT 462.470 10.240 548.570 115.400 ;
        RECT 552.470 10.240 638.570 115.400 ;
        RECT 642.470 10.240 728.570 115.400 ;
        RECT 732.470 10.240 818.570 115.400 ;
        RECT 822.470 3359.840 908.570 3467.145 ;
        RECT 822.470 2972.320 844.910 3359.840 ;
        RECT 848.810 3357.100 908.570 3359.840 ;
        RECT 912.470 3357.100 998.570 3467.145 ;
        RECT 1002.470 3357.100 1088.570 3467.145 ;
        RECT 1092.470 3357.100 1178.570 3467.145 ;
        RECT 1182.470 3357.100 1268.570 3467.145 ;
        RECT 1272.470 3357.100 1358.570 3467.145 ;
        RECT 1362.470 3362.560 1448.570 3467.145 ;
        RECT 1362.470 3357.100 1437.390 3362.560 ;
        RECT 848.810 2972.320 1437.390 3357.100 ;
        RECT 822.470 2940.400 1437.390 2972.320 ;
        RECT 822.470 557.100 908.570 2940.400 ;
        RECT 912.470 557.100 998.570 2940.400 ;
        RECT 1002.470 557.100 1088.570 2940.400 ;
        RECT 1092.470 557.100 1178.570 2940.400 ;
        RECT 1182.470 557.100 1268.570 2940.400 ;
        RECT 1272.470 557.100 1358.570 2940.400 ;
        RECT 1362.470 2936.960 1437.390 2940.400 ;
        RECT 1441.290 2936.960 1448.570 3362.560 ;
        RECT 1362.470 560.960 1448.570 2936.960 ;
        RECT 1362.470 557.100 1437.390 560.960 ;
        RECT 822.470 552.800 1437.390 557.100 ;
        RECT 822.470 138.080 844.910 552.800 ;
        RECT 848.810 140.400 1437.390 552.800 ;
        RECT 848.810 138.080 908.570 140.400 ;
        RECT 822.470 10.240 908.570 138.080 ;
        RECT 912.470 10.240 998.570 140.400 ;
        RECT 1002.470 10.240 1088.570 140.400 ;
        RECT 1092.470 10.240 1178.570 140.400 ;
        RECT 1182.470 10.240 1268.570 140.400 ;
        RECT 1272.470 10.240 1358.570 140.400 ;
        RECT 1362.470 135.360 1437.390 140.400 ;
        RECT 1441.290 135.360 1448.570 560.960 ;
        RECT 1362.470 10.240 1448.570 135.360 ;
        RECT 1452.470 3357.100 1538.570 3467.145 ;
        RECT 1542.470 3357.100 1628.570 3467.145 ;
        RECT 1632.470 3357.100 1718.570 3467.145 ;
        RECT 1722.470 3357.100 1808.570 3467.145 ;
        RECT 1812.470 3357.100 1898.570 3467.145 ;
        RECT 1902.470 3357.100 1988.570 3467.145 ;
        RECT 1452.470 2940.400 1988.570 3357.100 ;
        RECT 1452.470 557.100 1538.570 2940.400 ;
        RECT 1542.470 557.100 1628.570 2940.400 ;
        RECT 1632.470 557.100 1718.570 2940.400 ;
        RECT 1722.470 557.100 1808.570 2940.400 ;
        RECT 1812.470 557.100 1898.570 2940.400 ;
        RECT 1902.470 557.100 1988.570 2940.400 ;
        RECT 1452.470 140.400 1988.570 557.100 ;
        RECT 1452.470 10.240 1538.570 140.400 ;
        RECT 1542.470 10.240 1628.570 140.400 ;
        RECT 1632.470 10.240 1718.570 140.400 ;
        RECT 1722.470 10.240 1808.570 140.400 ;
        RECT 1812.470 10.240 1898.570 140.400 ;
        RECT 1902.470 10.240 1988.570 140.400 ;
        RECT 1992.470 10.240 2078.570 3467.145 ;
        RECT 2082.470 3411.140 2168.570 3467.145 ;
        RECT 2172.470 3411.140 2258.570 3467.145 ;
        RECT 2262.470 3411.140 2348.570 3467.145 ;
        RECT 2352.470 3411.140 2438.570 3467.145 ;
        RECT 2442.470 3411.140 2528.570 3467.145 ;
        RECT 2532.470 3411.140 2618.570 3467.145 ;
        RECT 2622.470 3411.140 2708.570 3467.145 ;
        RECT 2712.470 3411.140 2798.570 3467.145 ;
        RECT 2082.470 2975.400 2798.570 3411.140 ;
        RECT 2082.470 2851.140 2168.570 2975.400 ;
        RECT 2172.470 2851.140 2258.570 2975.400 ;
        RECT 2262.470 2851.140 2348.570 2975.400 ;
        RECT 2352.470 2851.140 2438.570 2975.400 ;
        RECT 2442.470 2851.140 2528.570 2975.400 ;
        RECT 2532.470 2851.140 2618.570 2975.400 ;
        RECT 2622.470 2851.140 2708.570 2975.400 ;
        RECT 2712.470 2851.140 2798.570 2975.400 ;
        RECT 2082.470 2415.400 2798.570 2851.140 ;
        RECT 2082.470 2256.140 2168.570 2415.400 ;
        RECT 2172.470 2256.140 2258.570 2415.400 ;
        RECT 2262.470 2256.140 2348.570 2415.400 ;
        RECT 2352.470 2256.140 2438.570 2415.400 ;
        RECT 2442.470 2256.140 2528.570 2415.400 ;
        RECT 2532.470 2256.140 2618.570 2415.400 ;
        RECT 2622.470 2256.140 2708.570 2415.400 ;
        RECT 2712.470 2256.140 2798.570 2415.400 ;
        RECT 2082.470 1820.400 2798.570 2256.140 ;
        RECT 2082.470 1696.140 2168.570 1820.400 ;
        RECT 2172.470 1696.140 2258.570 1820.400 ;
        RECT 2262.470 1696.140 2348.570 1820.400 ;
        RECT 2352.470 1696.140 2438.570 1820.400 ;
        RECT 2442.470 1696.140 2528.570 1820.400 ;
        RECT 2532.470 1696.140 2618.570 1820.400 ;
        RECT 2622.470 1696.140 2708.570 1820.400 ;
        RECT 2712.470 1696.140 2798.570 1820.400 ;
        RECT 2082.470 1260.400 2798.570 1696.140 ;
        RECT 2082.470 1116.140 2168.570 1260.400 ;
        RECT 2172.470 1116.140 2258.570 1260.400 ;
        RECT 2262.470 1116.140 2348.570 1260.400 ;
        RECT 2352.470 1116.140 2438.570 1260.400 ;
        RECT 2442.470 1116.140 2528.570 1260.400 ;
        RECT 2532.470 1116.140 2618.570 1260.400 ;
        RECT 2622.470 1116.140 2708.570 1260.400 ;
        RECT 2712.470 1116.140 2798.570 1260.400 ;
        RECT 2082.470 680.400 2798.570 1116.140 ;
        RECT 2082.470 551.140 2168.570 680.400 ;
        RECT 2172.470 551.140 2258.570 680.400 ;
        RECT 2262.470 551.140 2348.570 680.400 ;
        RECT 2352.470 551.140 2438.570 680.400 ;
        RECT 2442.470 551.140 2528.570 680.400 ;
        RECT 2532.470 551.140 2618.570 680.400 ;
        RECT 2622.470 551.140 2708.570 680.400 ;
        RECT 2712.470 551.140 2798.570 680.400 ;
        RECT 2082.470 115.400 2798.570 551.140 ;
        RECT 2082.470 10.240 2168.570 115.400 ;
        RECT 2172.470 10.240 2258.570 115.400 ;
        RECT 2262.470 10.240 2348.570 115.400 ;
        RECT 2352.470 10.240 2438.570 115.400 ;
        RECT 2442.470 10.240 2528.570 115.400 ;
        RECT 2532.470 10.240 2618.570 115.400 ;
        RECT 2622.470 10.240 2708.570 115.400 ;
        RECT 2712.470 10.240 2798.570 115.400 ;
        RECT 2802.470 10.240 2802.945 3467.145 ;
        RECT 53.655 6.975 2802.945 10.240 ;
  END
END Marmot
END LIBRARY

